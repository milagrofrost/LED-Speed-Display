PK   0jSU:e!��&  �>    cirkitFile.json�}�v�8��p�gn�iQ&�H0�������l:�餧�n�����,j()N&'�/�ϴ��H�� �V|w��N((��*� ��(>��y�������i6=z����2���~�����";�ȃ���ï��2v�]Ͳ��.�=���M��6uId�<�l'�	v������9z�����͑Ysl֜�5�f͙Ys�w5&1����f��C�P�~,�M8�c'�ar7��3c��5������	��m�0l� �6'�kG�O	#!�4��tm�v�{Xw)&�A̎E�ؔ%������!	)J|�P���T��� CcA�a{C�#ޣ:�C�,lF�g�$64�Q�=Dy���7隚t��lM�k#�bә�pj���3_A�:{BF7�6����!�B��	�a~_[J"�mE�r�P�����(LbT���$B!��7�:^bs)/��K�0
��� ��n�Z�Q׽�%v���M�
�C�����u�|z�k�0��Z�0j�Z��k!�Q��k!��������H�\����%�&v���[����?b���qL��;�P�B��88#N/�z&&�n�357̂�]k͂�@��8G}�Y��>�8��$�ڡ�P(�\��N$�s��1���Z=�EkUj��� EsUh��Qku�2����05%&��&]Yf�dҵѨ�LK7@5��ȶ`j�u��ռ?��j�jh5�Oui5�Oui��z3]:�@�RL+��0�5�m�q��I׽0׋��3}�G�I� Q`Գ��ݾYS/�1s_d�iV�=ktwϚF��z6�v��5sB��K�b+���}[=���I�>�;��Q�����A��A��A��A���J�R��B�u
�<��3!3z�
�IbBf��a ��A0r�!3�Ġ�0(�
ŉ�Q32��a�0�x�aP��A1V(8���b?t����� �@�A��d�Pb�aPL�A1�d�/�}�2 �|��P�%�?T�.{�}��].�O)��S����KW��v��>�.�����S7K��݌�v��&Ϸ�"�y���nJ{�,���@�;=�n�y *;��n�y *;#`�\�vϠ��1"�4�;���n���}��N^t���u����NE7[9 ����fw�N3!���N���B�&��b�ȃ�arϜ
�
�
�
��;o*|*�0��à_4~�0 F� a4��0 Fà�b<��x�aP��A1�x�aP��A1�d��B�aPL�A1�d��(�N�Sى��9����N�m����3��S���=s*;�����JE;�gNe�t��{�T��e����{�TvjZ;�gNe���N�S�<h'��R�N�Sٍ]��9���h'�̩��E;�gNe'/��=s*���3�R���.?/�}{�i���!�GG�i.��I��<��gy,��L6���e�"�� ��'~G.�m�8Ȍ!;�.4�c�c�4	�9h�|�M�<]|�������݀�L��p��sd��I�t !hFZw�H�L6Y�t�~%%MF�����	&�A#�3{�W�������������8�9�B�u ��	�����Z�m�����I2P�fQ����nK]�#L=��8�)�X2��\�:!F9a���l}�6��ЪMĭ�N��Ywݚ��ۈ���u�$�mơC������ۑKC�zC"��Z�����ۈ�����
B�7q<��PNQ?ȴZ�D�����u퓅L�+�����MV�f]��Q�ϱ49o�VG&�[3������i�:&��[���Y&'�|��S�,�}��ə�F{rL�6|e�H�f�����u͍�3~�P%�sq�}�y0������;�)� �i2�}�cH�qu0t����D��E�[��f��9uŁ��3fyu�}���7ׂa�ߜ�e� ��0��DM
F{�w�p2�=�d����;�]�û���~t�}%�������l�5�]`��N�>� �3|:y{�&��t-7Q�S� 2�~8�U�]y�<|GU>���8y+�x�|k�盿c��ph�O�-��>����!�ߞ_�}�o菍�,�,��l����$�D�J0����C�0�L���D���3�rp�]�J�����qv̊�m���%�n�%��;<)��	���H�;����Ht;kU��t�
��i{dt�}M�*8Hx�C��_uk��f5db�2x���u{�4�m_�Ep��_��n@�{���pK� ���{Â<^���1���Yu��<Cq�Ʀ'(��@ư=6lO�S��̰�<U�i�1	*=Cv�a{�NΦ<z����F�M��V>��E��E��U�!0E�:����p�&=�g`�(FF�������Ŧ�Ŧ�U� ���['Fy�J6qU��=k{��[�25�p�&�&��&Ʊ�)��)���/&�(&[|���&�6��OAl�Iz�lrg��j�0�{d�}4b����F�����e��a�-r=�:�S�d�}|b�������B�@��� I�d��#�>b�E�g��>k�E�/�{�b�\ϼ�}�b��j��h�~���>kѤ��%����-C���A�zn@����>����"�3�h���"��B�cl���*ڧ2������3�E����u�P��tpg�}�wH��&��2���2ݨ[�o@K��<&mBBE��7KIJ$J}K�+Y�O�Z5Y�)Fyr5; Y�H�PYf�h�X����z�e�V�X�cC=�'�Q��D� ��- �yW�P�{p�X'�m�*������� u|h���h��it���@��c�0�FO�d�l�3,�/�v@�D�ؗR��1�8��k; K��"�ǈ�n�P�w����c����{�ؾ� �'벐FI5#���Ďq���P":�$@��E� �(���� {0~��A�;�<�1\V�L ;�K<�u����8�A�� !G��HQ���Q�1;�ePCCЩ�>�W�]n�Y�P�rPAH��fQ$p�!�;�%�h8ȓ�`4����,aN�rD>���@�nAh�T�(Cq�5	A��1(�A*����]
�7Lp(k��[�m*ҷ��[Ε�|��0'#n��nn�ƍI�e�t6z��!A�G����I<k�Q`c ���'MmF������D��h�ϣ�L��x�#�6wnLO��\�t3s���6� ����5B739tjsI�c܇8j3'���ANi�̮pc|p�fr�dN0=�i3g��N��Fn����ͅ�J�$�DƜ-$s����V��)���"�,r7�pY�7�����,�e�,Be�,"e�,��"o���E|�UCF�cF+>6Aՠ��Q�$��U�F��F�fЦjP%� =��y�� � ��y%��$�/�BR�~�bX���rz���8��c��s�����R�?�|"�t����m�'��t���4@��G1��s�A����8����a�x��Ak����S�������$%����}���ς�\�}U���l&�E*dI~8���4�B�Ǟ�;��ݐ�P�F�"�F4!$J\0/�eQ��q�""�H��_�t��Q�F+E5:��X
N����4�&�d��ͼ1���\�|��)n Z�`oL�r��jª�l�*R��9*�!Rާ���[����v�򾏻�#�ՠ� a�S@`�5�a�^O�k������E�&�g�&˒MM��,J65Y���dqS���M��,�oj����ɒ�MM���,�&��MM���,65Ylj��&e��1��ˈ7J�I,����G��J�?z��h�Q,���G��Gi��`9����QX�Sqo�Bl{��4�I����<�d�������(�r�K�q)��*�W1Ī�H�D ��h+��� �f�z��M88�س�L��8�<q)�j�b:[.j�EHp䇞���Ա�DؾG�B'	y1����oB��dm��k#yz�N�e	94��[v����&�	"�ļ!��A�g��31�%q}��V��>��
���I���l.��$������e,J�',�(A!�w���ϳ`
v���^�!�������p�(����W,�%gY��9�s1��e�Fh�{��t":�4�VuH�1���	%Xx�(��4�P�i���R� �r@�A���W�k;��0J`�C� E(�&a�G�0�3�
.</�Ŗ�ƽ�r�VS8���A6��{X,��,#�j��q�C**~�?:����S������0�-Ϟ��+�F��ϟY�h9�B�PKU|{�έY�]����K ���T�E�f9�M 6C� �ޔ��t>�_�+Es��,`(�?���[�u�e��?��k���6�r�H�^\���hͭt
-�_�q�b0���ZV��0r+�B�7��9p���Ȣ�e@�"]�7�v2D��25l��������a��=Ǻ�L�KY&�e3
�Eb]��5ϒ�u������b9w�3�DA<!�PU��?r ;����P�2�B�Rc}j��g� c�W��a��|.[�K��*!Jj��0��l�.+�U�������/���Bk9��%�h�V�c����R�ŕ_p8ɲي�x���0J9cY��+��/K�J+I>	d����"����Ě�a�_�v���`j��
^N&P?���ŋg�WU��ip!� I�0ϖ0za=��^-�B�Kή/��Up�F�e0�*5��S��tM���޿�fj|)�OO����8�襋���!�Y��(&���R(�����s�'�<sF�)�ͱ�Z_����T��K�/�n���ٗ� l�ؤ��Be\H^�@r��_�O����j>�:�˟d�b��j�?�	�1���������KA�U�uz��eG�)��YQ|�X��OOAx˫q9����tq��2ab+=���]��/�ifϗѥ-'��4|f���:P��|&�~���Oi���� u�9���C@W`����	�z�Y�n:���H<S��{��:L�*�X�;�~)�4Y��*�'"$�$��*��td=�|Y/� >}�fd� �Q��n�� �Jq֡Y��08W�G���GPY:N�m1��y�C�H*	:P�*_.�r~���NS��Bo�����U��#�E�eu���RSݪ$�Ӌ����z��h�^	iT�-�Q�QZNWo���VY �F�<��lU���M����7�%����_�|�?+�:%��j�ra�v��YYm�-�G7��}�V��/�9LH`��%���G��e�[�b���l���-m	T�U�
��=���WO���}��s�����	,�A�K�u/��A�0�p�Xd���Υ���_�j�CL)fވ.�4p���R�0E?R?�/ �<�����mk��9�����7,�>��|uF����������͍{p�qw�{���W�l�+n��5�C�{�K?����Q=Zo�S�]�4���ߑ�g#�����β�I5�ZE%�jy�W��rh�U� ��2BR3T�|^Z��R��:vl� ��*}%=]��*����"
s+)��c,�Fu��\<>�%O�%�m��d\�� �W�K+*���5����+֛A\�fiJ��DEv�"XN ��/�*��L��L�y¨d9Q�@:M��5����U�Tj���&.�l�X�斜a2��T�N��粋8��#I�O/D�ɨ�2��Tw�&S���֒�&قH�Z7�{�
����cխ�am���S��k8+�TAZ�
�`�ʿ�f=�B�96�T�Q�)VhE�
�XY'X.�J&�-)��k�������p��ԣZg0��"�䔼+2��oD���&��dz���<��A�����GŠ®���b�j���RD%�gg
[�\�-�xGV�DcX*=�]�\��=*(?���eL9>?;S$d��CKI�����n� ��\rq^&�gEX�RĩRD] ���+��=�r��O��nH���%���!�r.�a9�5V[�J��'���ã�&O����J��ג��Q��`�W�_W��P���_(�����fy�m5M)�[���z��U:��s�k��?5c�5W�@�����Y-��eP3���◿�x�A*>u���t`�T�֋)L�$��z�qK)���q%=���k���b�F9���G�� �)��S���ɢ\������^�DU¥t������\Nmr��|�^B�].qv=-������XΚ�E�������Kшހ笭$d���lx">��u�l�Nք"��y�T$��G����i���
�r�|�q�����~{~��˗������x}d���-�X��Z)n����N��bD�Ry��-�K�8K�o��ݒ�ɨ�JX;���W�<�d��;�R�J���tz�ÎS2)9T����r������
�-po��T�o�hu�.��lM�֎n=�r��B�����zY��r��'��HE�J����
V���UmN�:-&#E	�wk+����=y���7E-o�^�.���+Fs�� ���+zL��޶�ھ��c5��2�t��Ic*��l��>	J�|���G�[Ū���^@��:�-K����!:n�s>�ș�F��R������Z`LV���_N��Z}��n�}�j�n�3��Q���o��1L���co�o�ڻE�0w��@�?���;'�J��u0���̔����R���M�k��%����:�njǤӎ�V;&5;n����8[M���")�b;�UUx�e�Wi�^��DX�y3��uۦ�h6��E�^�q�>x�`�j��.3(!mԩ(�|��i��D�<�@��kQm0]���qv���b�k�[Xn�0W�wh��H��"]qw���5�X�V����fB�O��d��ht(�+u�v`�����vA�K��Z��g����5�N6�Ѕ���Ю���3����z?p������z�v��v���s�ѩ�5:�kt�����蜝���wt��٬�?�ұ��Go}Sx}��a�;��[���/zT�v*Mp�R!۩4A�v�2��J-�^�fr��r������ |���L�d���E��uK=�l�I�E�:�Fٕ|4��j���v�8��d�ڟ�a=�l�z��#Ŀ��I�S��*-r������O�G��M�h�b}���Ȇ?�����A}Du�+���l\3��i��x!�����Uv��oݾ;��o�Bmy�j2�;m~��pFVo�V����T+�Tr)���#�V�eo��|/w�қ��Hz�X��s����bP.y�̈́c}�`�����k��G�5�Wֳ�XUK4�6ht�\l�G���f�U���\@��T�|�T�㶎����Ȭ9��|-C�����h�jb)�K��21T�{#&�&�b+ⷑ3:*6���ot��om�F��c��=J�)��8��!�y����9�6ڹgc6f���h��Wm�e�1�����=�>%"�o��n�4���(����1�����=�Z'!h졗{��SV����1�ڛ�˂�VmT��Ucs	��ec1�1c߁;E������)b�1&D���\�Y�bW�^��m�i�����ky�د�p�?��N���Nfԫvd��qG�"��0n���D"!��>s@d1ŝ q\�I[dZ�_h���m�Xm!gNqe>t��SxY��PØǝ\*�]���v��K"����c�:�C.h�}�+t���]���ۆ��)Lԡ͗�h�@GA�W�kA�Z�o��xT�t�7"�c��s]�NsO`b{!�&�� id�0񜄸��E[�Z��h(��V����;&͒��&r9�M�ӂw�K���2��q����Vit�e�Iԫ��i��������o�z��(�����4q�ڦ�or������Ć����H�8�6�����,ҭ9Z�Z3��,�:������j�-g���/u��_�O���=�:��.���Y��N�'�Z�o�]��e�I:b#W��V\�1G�� ��	M�5g3y�1y C@l�
��̄HB���I��@@1�˷���=>�}�i3g�4��7Ƨ֡R:�'�Hw���a�J]�a����~+������Z�i�~e( _v���=`�+`������`��<�Z��cgS�j����u!�|�����`	����Ή��$TAR2�b\^�� �I�&�"k��mUc-�k���_�i�8\��C��l���K���֪�ڝ�y`ǚ�Nm���I:{Z��q�F��˳Uߪp�ǋ<[N��$�kL��i�Y��D��>�u�׳ j�����֪���<����ui��"0��u�Mo��N���Q��X/�gO�% =�^��m�5-�c�R�0�3��`��w��'�e�z3׭�)�-� ��������Tpb�(	J<;I�L��Q�m����=Й|e}^{e]މ����*�,���o}��hګ���򉖭^/?�7�?�F���kX#��c�3�sq������_�z�v�u��+����f�ʺ�\�����G�\��H���/����eֲ����	u�OG>���e��.��ek�R~-; k>�O�?C��to���yHˤ.s�>���)�hL(�b�0��cKk}�Z����x>��rZ�r�<�7�{S=��b����_����3�u!>f�v865U��r�w3U�ܛ꽩�Tm�KB[�qαG��R���`)�qߥ����]�;h�e������g���yo�]�"gL��`x1v؈!:��ܖD�aDL�R�+Tw�.���m��g�cJ��&IBG���R�g��j�����v�l�57�O�,?^�P��]����v�a~��1��0�ّ3�.%�����V��)�!�,��x�N����{{<�*��r�(�Hr]f�F��5��A�#gg|t>[z��xc��"�-�;�`1L�����r�#`�h��(b����|M-R����	�A��2xa��T�Q�Q��G6�t�<����i�����ѭJf��K!�×7	�����}n��R'"���R�OV�:��b�����d���~�� 4��z��#�?������Y:-�r�o_@��[Ii~CY�ʃ�7C���Ȟ:q�,X\*b_�����h��3YP��?�w���WUWc��r��0��6^RY�����X����},5�Q��C���3}`���P�(���[�5dPօ�v5�vVk���W�m@q h�#�]���j�>4���.l��ޞ�إ'}�c��V�M$�1`�}���c� �Y	y�+�q�oF>�3K�����%��);���^ҍu>�����}F}ֆ2�ŋ�O����@�{�p�*��F��*���.U��ݞ�����:��pQsq�Y�O��8k��u���Z��������/֊��S���V%}g=�����V(Lָ��ރ�}-���yԙf�}�pm���}�g�ZR:'�f�{�ZysA���j�c�:j�7�u��ʛ�y�l8����ao��.M���y�B�_K7��T�s�ΐ�p���kCaý4PSM��M��wS��<�e�{�{����=��W�ͤZ�.թ��Wӝ�_���=f�=XJ�7� �V��8�u�j��u���ˀ=��kCE�7�:F:���QȚ�n%���TO�Z��=V{����=��S�̩��n�VOb����!���������m���F���w�=�=iڰf5����Ժ������������A��x�>��hw�ػA��èc�^W8��p!��x��o���o���톺'�a�V��3e�R�Z�tݐ�QL�C��"�b�C��&�hw��ݿ�.���a�K--�4�D��E� G=QNcѭF��_�f,�S�Ar�n:��N~�CS�Ts�#�����`�$�z�Ws9�ߎ��?PK   �dSUv_Xh   t   /   images/0cd87e23-7b82-4f28-8831-3bf70f36678e.png��s���b``���p	Ҍ ��$Uo��q��ܝo�ԩr8<"���A��a�	� s�O�������>�ry�8�T�IN ��=�/)�<]�\�9%4 PK   �]SUs� ^  7_  /   images/12e44cfc-662f-4e22-b257-55fcd330266b.jpg��P\A�6��נ��[�ఋ/�{pY�5��������!��$����u��n����{�S3����:�z^�_� x`9� ��� ��D����DU�$�O  ���  sps��K����{�o05su���g�~�?= 0����?������x�����s�Ϥ�?Nd�������ͣ��]��<�g��o���nNn����9������0{w���7�����ƿQ�_��  y��������|:  �w  R��>e  �_ ����1��7 h�r2u1�_"��� �. �u �i  S�����������U����,�I@ ����| p��� i 
222ʿ�:�?�baa���% ����'$�$%$"'��'�%#�����!$�c��f�������K�P�p��q������?����A�GB� �# �#���  @C@�oYF@DB��I �?�!޿WD$$4TttLtd��h�(���hܒ��Dt�A	�3���<��$R�O߷�Hy������Ps�/}�2�!Ʌ;�4,\0�jj�4��3O� @@�: "��"��S��H(hH�(������P�?�y �	�ļR$A���5��^W o����G�|��2��ӷ������f�>�A����O�'=���D�L���jI���Fvz�K�h��O�u�m�͹,����u^ٰ`�h�)��`JqA1B���=�H�ζ[�k�IӺ�c�ص`�J�͹w���j�L�N�TK�٪��|�|;�b�GA����/y�
mT�q,#���%'��\�?�|�m�e�(��`|�`?s�*pIP�6�FE��2~���U���.��$�'f�WW4D������F�>��\�qv~�3(��p�E��w|�':�j��l^\�r�v&f���C?ki�R嬂OQy���}������%�gݒ�̐�5j�
�y�:4�aV���U�]Y�����m���c ��4]�R�6`���B9�f �$��(G��?�iwk���y]�%�݊F��+$��6J���fE��х5��}SZ"TRA��W���c[{�9����@@ߟ��ݦo�^��aӓ3�
�]��^�(S�<����CYĆV�>�>,�� 6!&c�y}����I~�?�`E�4  j��%8tVW�|#Zް�x��[�v���M����7�o+ʘ������c����	u@��w�D�
ǎ�h`s= 1�	���t���1&����M!��[i�	��D��Ζt��cr��u��>/_iz���s(�o�A�|w�b7wڐ��.��~>t槤ģY�_Z�1��|[s����O��6�Y��8�����������Qn~�˚�FO��_rf֝Y���|��ǽ��<}Ў]bxIJ]�^�Y(Є��o�1��Q����U8}s��T3��.��^Nn�W �f�[���*c��,r����E�\��u�sg3��Ƶ�^�+�����`�i_o��ҪWGj,]�-=�e6��+U2��3!4��N�h.��=l8�Vc�T�G����-�R�h���j�/���'�o�$	�U��|nG{�)Xm}t���ā�"�����%%-���ze�<���I�S�(�R4s�w���m+(�׵�wW.��8��ey�<AX�@����v��m��h�x�gy}���f�%��0�t�������t�s�z�B����T�n���ڳ��H��^��W�01��Cvd���cП+����h�t=as��,�a��Z�;�-%k�w,�����1�&3�f�	���u�c����Dk���X�v��L+�S�^�2̲&�WSgnT**�(����䏁��Jm���]Hܛi����jD��J��eX�߳�����Z�ۜ0����g'�룮���NL<Cq�⁼�K_��#���)��6=G��_R;����36o��M��ܙ�����+d)�?�>B�w�:i��Q�=ZAwL��&b��!���
�c�:il������_S�;����A�Am���~Cɐ������S��[����S|4g������2�rm���-[3��]�yK�plR��z�%�@�,����@�Y�� � �h�W9�^��+i|��!
ŧ�p��|Ǜ��,�3�����ͳ�%W�����O�dV�hc�7�Iw�B1궟���=�Qx�L��.\gҫ)���Y7Dڗ�~G$Yʉ��d�C�x�i�2k���)x_�^{�=�j9�V���D��G^-n�89R^2}hYL �����W����ɝ�"��{L���m�Y?�?G�zSf���yw��U���7+���o��%y���0��=�Nړ�
Ot��* �H�o�u��]��"r��]U���S)&�E��7d/��t�<���Q�9p�q^0�i��L���*�OK��+���<�3Z�[U�����S���Z�rn
�H�>�#ײ(�k)�+k���`u�I�#�N���H��g�wU����t�CSӮۥ`�����{���bP����� ��a���cUɹB���>
6�F��X�C���QF.�<��6�u��4���*nw�1�� ����EAֽ��-W�|t煉�N05��a��$�< �T�!C�qG9t��Mj�/��Lǅ]kM���v��jf���c�I"��]��G�\�o|�g��)��l!��UHM�T[:k[�o�'T�e����P���n�J)�5B]+$��U=�dQe@�\��A)�A�mm��%�f�mC,Gn>������Q��%���0\��;fj��O'��J�7�|��z|9�)i��E-��L��D�x�N��gg:�(.��K�_�_��`����^�3
���@x��~Q6dze4����
jJɼ��I�)�ƣ"k�A����բ���`��	p�:���U�9c]b���0D��h��1��ؒr�X%��a�B�j���."?G�=Vd+V��IC&���}��7$H�	]J)���[9S���ڂo��ۆ��@��^�]�|�},�����PR�>-�~�`��_�m��zZX��tn�%��[@��l��S�.�3{6�F�tP����*9�bh���s���z� �tV�j�-����4d���,W��S�C	.�Ԟa�j��so^��%��tJ��<,��qxs9#~'��$Lݡ�TFE����ۓa"�k.:�<��u���W�G�m�g�{��8�b(;o�J֔���5�3�6����Od�`g�ޔdh�I̚�(O.�kU�X�����ص�F�y^�����$:��LL�25��^p�i��/�4d�[7���� ��h�Z�&�{Y�^b�z�JC�6��ǞW ��s/̽ěX���${�@9ߧ��W��*�,h$�@y�B<j�]��8�N�߅��7�34:���ᦣ"�\<M�7�� ��t�+��R=�*W�c=G�1����)�_�(%�i6g�������m���`4��#��nP����s�$TJ��#d�Ŗ
�#�R<��sẼ���|w^b�v�p�u�iFF!8ȸ��y>{z} Z��D��Ǫ��fb͵�N{IउB��WW�<C�A������k�ZA�V�܄�7[���0d�! �˪�4iyg�E*�� '�Z�t�ϡ�|A�\UcY8�P�E������0}ٗPm��)�|w~�|8�ǂ��U���;V,����ӇV Q3zC���*ב!"�0�lBiRߍ}ɰ�b�.0T����+�XF�� }{�*�ѕ=T�S�2i�ݻ[���]S�Zy�3|s@N��� ��S��}L'�G���E�D0u)��	�;\B0e��	�Z�Brq}��ZU#P��ѴU�pp�U�/��۾�y��-\.�y����Q�ʪ9�V�����
��<�r���3y�z_O����+`���z&~�Y)���<q�J��%����̐��%�N���?H��Mֻmh.��=qy���f��Cah�|;]�+ 3.�-aJ�+��|�­��VR\:��Y��'!	�W��x#�>�«l�0q��_.A3� �BC�[��A�4�p�D[vj��%Ø���}�@1��d�+X�Ld�y�%�O�dM��"��W�6�aB�A����Y���<�n03d�kx�Y�,!I6+4��&���e�ʺ�c�}�����8Tx�"=29��h	b��'��A���c8������Yd�ط�7}�Ѯ$�^.֌�%�MP��@���r�;���=;���y������u����?����=���c<&�8�A��zb���X
�=�US
\ͺyZ��6.�-�;�����2�\�l�͋�����?u5��]�&)��e��,�ŧ�S�2��)����m���Ŷ�r*U4m����ӌ2Yl<hM*��/ď�<��K���X���()Q��Cђ�֣�6��%����~����ݾ)*�g��J�X��%�%�}$#�0�����Ǥ�>ja&��.�Ԯ��;����������2c�=�ڟ�yս�Q������Y��,<�]��	��:5�ڻ�Y�e�N甖0�<�q�o$�����k�*�&(D�p�V� #�>��b��b����N��F�E�-�"FXչ�2�ۿ)������xk;"��q���|�|}�Eƹ!60.�PF}�~p����ª���($)�@,/��.gg(=Qp_�$WMb�Ё3D��<�����읬��G��&�k��<j�}��5�S=�S_���R�9�Y�z��#<.'�O�TŶn��b��A<V�E#;��)jF��\,��og%�Mr,�9J^��:Ȼ�<L�7D���� z���
w�]Ԋ��?
��v��ɡN�Jj�1��b���3�c��_����EF%Gv��+��vG4���\�AOYT(�(E�[$Vy��*�gI�����ߩp��KHM�z��6=�t7a���p�.P��ꎭ���+��=�\4�	(�hU#�B4܎5�*"���8�r���o���ee�橲y�-,��>�,�}Vwz���y�b<�-Tƶ����2��á8F�/t6�����Jx���0Er�Q��*�ש�QIg���3�v�WDt-&�]=��:�
xCʨ���)>�+�vR�s���%����mlܼ��lˍ����z:Mt�)%�I�� ��O2��5&�(���!��W�r���Ƶ��D�zvO�ϤB6�x�EkD:Ì�9����XynY���(�V���ƉR�.:�5*���%�,9$�l��*E����g����H�lC����giu��ʨ�&���~���+`Y��9���@��_�i7�横u�]۵���T`�!;��R}�����qfI��@d1�]���G%�W��~2P�'m&��oLb5�W�/P2�5���u��]��.H��c9�q�-AEo|cm@ IR��/��\��)v�&'g�)q��J���\�c:G�x	�y���g�C��I��Ͼ�.M�Us����V4~v�d�+3:2����^���Y��nV$���:��˅k�n��Ө�ڜa�<�&����h�Y���at��|_��a�	6��$�z��Vd�������i��V<N9� QU�%�<RWOY`'{������@J	���7���'e�����\�$'jf��Ń��ȧ��2��4��­[�@K�Pᘤ��xe�$g�Cv �h�×V.&H��Ag�i�w�O*Yr<��}L\c��*6���Ǡ�k���7�8����/6�������E�bk'�L�,j�� �skL1l�}�NE��<$&��5x� �/�-�F���%�E!�N�R[Dy	�M|>��Z����TD������X?�1��G"�]t�R�
k��ԩ�rJg��MDވ����^�|-�C��Xa��K���F娥����aB�:��G�CJ)-��a�d��y�Q][���^�>�&z$�LGJ�+c,`��jZ�S�IV�dk+���qR�N�%�Jp;�IzQ�y�=J
��a��R�.�a@���$����)����1��Z��Y��|h��f��L��g�6��Mg#g�{�pX�I�G�)�1;$�hP;ɿ�$Z�r�=�J#���m����k��YTS���g#�Vťd�YP��a[�2�K���8@]Q ��؎�f
��kL
 �X�A��G���Z�Khb�V-��w`�A���G��+dt����m��b�sV���"�/��1��G���Y�:���*������1j�3�a!ԒI?�xnr�2����;Q�Y�~�����_�=�E;h�� ��>`�kF<�*�Ӎ���	K�E�n��"�䰤}���RS���+?�
������K~�]�����B�Sސ��+�3�h�7ӊ��@�`���x�\Q<KO��"6��y*������vds�/�� �ި]�:��}���EH5���d�ÎV#���ԭ��a�QZ�h�.�j+M��8T��"�I��S9~�F��6n��N�\�^��+]>0�2�f��U��	圐/��t�$�-1�����uC�V���B/ּ�-v��p�g,n����W6��'&�z�v?�#;ѯB�LBK�g�Xg��$yș5&�4��AE��@A`Nnt>8��iA�X߰�k�Ƹ���6b{i9m�I�$2	��ni�ôI���ڽ���;�wqtg}�Ҭ������8(&؅$���x��F�B�]>��n�8c��+Y�/���hњ)|Ia�[�r���ع200�	/��������j~����vF����,���Q�R�	���6��f}u�u�Yb��]X�+�-�y�[Q� ��Ԗ��ΏlBn�����h��_��{��6W�JT*�lN��	�m�~[f�m����B�b�ov���CZOھ�t-���|c49*�2�~t���#���nS���S�Z�Q��m=�jG���d�fgԄ���Ǉ&��F�⯇��T�����J"��ڲ��ڬ=�T+�M �E�R��6�7GM����VI��2mA�xD��Iѵ��ጝN�Gn%r� ��.��i��S���ӡ�ʕTE����aDc��#"џ ��[���T��a�Es$�{����V=�}�WG��ך��u�'R����S-��5�~(7K����#*�R9�@���g��|�r����s'ٰ��5'�YE�� n]<��Uڶ�?('S�ʢ�n�!��ۻ�n���/�ө����F��e�Ms%Q����E˞�v��������\F��>=��7��y@�Bkȿ�J-.�
3����)첈d��=�.�Ȃ8���؎h�=YV(����9y�������g�W�))�
��c@a��1�Q����8L�B��9�Jb�^���_��:�/�۰z!�gF��^|���Nn�I�Z��ʨ�5���o�4�s'�2�JF���{��P��B)�uf�X�
^9jT��H)��*�V������cO	'oGl�Z����~�M�&x}�Od����*c:!d��晡�d*��do?��	R԰����ȅL��s)�,��3m4(F�M�.m���[y	of�]���2���Xˢ�	?7e���՞n�i*�u̿��0�Wbd��t�����k��t�U\%�g+W쭔�W�i%���bB�Z�M�tn�����߃Ξ�+o��T�+�k6Q!�� w��,�nQGZ�ғh����V`�\�"*�k�@�Q32����!,��6ʨ[�H�z�*g��ӵ5��_����[V�>!y����z)6E��ĥ,�y�&�w�G,�x��9��r���`N"C~x�u��ȹ�NR��<���%Cg�$Oh�EO�u�{5�T��Ib�h%khN-]�fz��U����>�U�)IU�V�N?�?	����Pr��)"�JAa猖��@�K�p��L�#*!�]u��.|���lri �ȟ��vsǜ�8P��|'Z\V���S�F��,��Z���B��m�T� ���Ʌ�B4�h�`Rx\P�B��t%�L���	)���^�$��LNz{��\&�~� ��Qm�f����ecE������+߶��fF��T U��D"��pQ���]�cC���'����#��J��F�B��9yU��>�.�G�w��Y�����zBkf��m_
��Q��$
�l��*<���w�y�r.�3�̬�L���9�'!q-����GZ�]�6/���왯��^N��^�[�I܅��/H��I�~��+��x�oa�rh-��� �O���J�_������>�ϰt{NS�s�l+������3a�� Z��������:%�.F>��a��r�c�	�Ád��ݣ�,�p4u�R��-�{1�4��9�)r��׀�k��7�w�0��B���(���&���{7u���r��yh�����V���;��E��z}�u�'�'��Xc<�+K�����F|�X���g�f��Ko4뽃�E��U�GV9�p��m^��#/��cX �<����E��]Ї��>&A{~�j��Hf��;m_| L���LH�|;4wootҧ��B�����~�_a�9��Ez��� ��#����/(�E����&���5�Ax$���R�n(�Q��X�Z~��Y4�֔��h�:��X�0��>�W�,��QK)�#£ �R�waN�29����S��m<��?I./�#�ZeU�UT�6�	B��MI��3��n"������N�A�����;�wo�o0��;Q%��Y=��6�!�5�h�L�U�g������o\\����e��c�~'�K�?�>�N�!'��j�WLSX��A.8�ڊ��>P={������[afHG����Nf��j�����^������X2��z����R����,������I�)wߜ�Q��Y��u����1I��;r���R;�	ܱ��O���k�fQ�N)AwMy�T��W���ԌE����u�c��ύNIn!��������
��"��?��8�m����}�گI������jU��\CCtFU���w�j��&�1�p1`C燱B'L��kNt�7٬�����ښ��5*:��Pڝ��6Y�Z��w�󫒜+4������UO�ȐC6^������<�1�����(��r͟�����u�k��agK:_���E����U��m.�=��'p�Ul����2�k�-�Nc~�v��˰���#��� ������W�zI����Y�p��˗7�dY6󱯀!��Ę�C��s�~��u=�0�������ʿ�05�ܿ�������ۗC�~�w����y�Z�\]�XB�l�V��މ�� ����̾���5�%�z���̠�� �
(����AE�6sOb�1���gY~�MyC��a�M]����9G��,��7{Y���$���c3��_3�֠�>�W�y�l	��ƫ��A�WN3e��<~�sw7
ʌ�>uG׋G#c�:���V�?:�4�i>74�T8�SkD�p<����-hq��]�5�޶7V0���g�R��m,T{�i�P'���W���9HT����7[���&k���<�y�Ei���S�X���o�0��p뒨�E�55�T�,��x��;��r�ъ*�-澵�5��l��~�e�Z��Q�W�OM�Z�*Ox���������]흫��4��BMo7G���1N���GJ���9����S6v�֌����A�o?1�7�^�,�=7��8���[�S�w4X8���u~p���%����%35��yI%y'��,K��G�cq|%<��h��	�x�1���������|AW�Jh{��U��C�=<G��H�Kih�ɿ,ФW��rY<Z�pe�9��2��S��J�UH!g_��b�Σ��\8;m��~��"I2~H���M�c�|\�r�§��s�����2h�)*�VגT�2W��s)ā�}��C������>��9�z���PW�$7��D!Gԗ���\uƯV?��,��C�SG�vFheʼB�nN�x�����υ��:�3�f-���A w�=�y�Z_�m�;=��&<a7�]����3�ʘ����J��t)�Z��QlU�gÅ�9~�ѱ�"[!��|ݘ9�h{��k�e�g!�vs���h<�ޜ�ߏs�1�T.�����c�����C��<5���`g_�F�?g�ι|���$^�������d�Z�6s��x|�l�&|"����<�էT�#K�� ~�Ce��~p}Y����-+�I���O�l=;'ȗ��R���,͡?:�0˧�^�W�Ɩ	bSSecH
>�$�K�>����nf�fc�-��8�c�^7^B��������. :r����A�q.�*���)>>��秒Rm��3�$*�41z��8)�;d�����-e����0)�$��g�s�Κ
�L� ���+�ebA�T(�K9��HiZs�s��0��
l�$��RF���M\������u�#�+?b�B���cNV��c�c���aOgpp�������끿Ѐı;�Kϡ�zٗgG�g�rO��Sj��X����(����k��?1:F��5��$���7e;t^��c�o�O=�ǯC�v�؜�g�/�t�k��a%@�Sݛ��&���W e���4>����x�uo9���:���W@�o�Kܣ;[��yse^>�;���	zjٯ��z���+2r�/Ex�����GE',߾j��-wt�W���ZŹP�+L#P��(�Z�ќט�9_��:��9�n��=��-K��-���P"n7�[�v���^�$�ٲ�hۦ�
���k��G�٢G���U�D�:b�!!CW��<A_�_JȽ� m�>��9>�r�x�`eL�^��붩��؂�-�-�y,��e߂���%W�i���u l6�?� ��*�N�@����9���5D����q���u�^��*Kf�<jNI����Z�,Z&2��x<��co��C�����6�d������NT��,�~jD���r97��Q
���2G�F~�̰��״��V�T;a�L���x�9N?{)'U��-UNlz���b�H�M���(�W���&2��D���-O��\�6����ۼ�E���~|�6����������7�b�w�z��l��� ����#L_9�ѵs��o�G��I��IRE����]�
^Yb���k�(gK�>���POX�}�g�y+fML��eZ�V@�G�A�G#n����H��%�b��l:Yx�*
�+�}C(F��޽A�I�7�}��W�ѣ��#P�{{{D�tQ�;`�?�t�?��!ιCf>� l��ѻ!/�4A���+y�a�F[:����h|+~&���BRW���8����;�i�������ϞN�)�������]ٵ��	.s��9�͠.���3{e'�MJ�&$B��r�C���H�9�-F���ً��ax�[̌f:$�+섃���i$%n��7�~ڀ���n�71�QSϕ55-��45$���[#�<)V��t��f��#���[��1�n�׉�Cg>l��6��t2b��,�a^g�k�!�O�Sh�ɒ���cj�MW8c����JYz�7Z��#!Yڤ�A		��-�3J�Hw1�Gf(���<��]���,n���-/9�Yz��/x��t�D�q�� =��S_%��ME-�P#u�c!V�d�iw�XiqX;���˛S˽	�@��NB�YU�V��ёt�U6ZUO��B9��J]�� �����9��ު'$@}��t���c����2J���Oi�]pc��¹�Z�ϑrX��a�}���1��m9 � U۫��
�[��1*�Il;���3�&�k�l_"B�_.?zs3��>1
�{���i%z�g�����+dE�H�#cQh��D�	kr��g'�.�]`����H�w�we���ұ��ۿˍe�q?�C�R��Ͽ0�D��@M�8�J_s�bL���b�&#燐�uI��K4V
bچЃUS��z��u\����fN�rEB��K֬����Fzjr��C�ڷ��%���5ר��/v=ū�ʟ�r?��%�~�0|}_zv+�0`�b�.Qߛ� %�����LOR�F��x=1g�$���V�	WH6�BGw'�]
)���bZ���ߤ�ܟ���x�t=���4�%�"���MT���5��,T˂X��v�aǫ`���E ���!�VD���L%�J`t`{$U�|�h��U*�GMO��\/�t�<}��N���V@]�&q»��*��d\K��ۋR�ǎk팎X��6� ���~9���|�� 9�6�Y���|h��o�1Q���횣��t�0 h� �+97N8}���'3:���N���S���
"9���	K�c���_��f�P�c�F_i�u�ޞ�ux\��y�۶|`��Cf0:̈��<�e_�,Rvxd�?z���Y-�Pu�_$/�(엽����]pO���B~����6dkZr��r\?�\q�,��p��ۂ�p=����H���Djfٲ���˄֪.nH7��i�-Wa@)���i�CL}��&��*iôV#�mQ�ѡw�y�wUt�
��7h�%w��)�ܛ�)��J=���i(��v�JQ��RޒO�ŕ66���ť��Qi��aD_IQh�Y�|�L�5�fY�U��E8%�%��;ֽb%(+6�8Վ�!V����z��
���ݒ�v��`�O䟒�+l�la�F��A8+`��~�㻇ؿ�������߱�i�J�Q���|�� W;��gTy���<?�x��S��2���E� �K<M�O�aU, {�wyQ�����ʂ��=ᇾ�L?��e��q�bTy.�;A���+FR��o�ӎ�h�+�n����z���pGE��(Rm$�!!!��O!��o�Ұ�x?�9:�����'�À��uzҋ�6���3�ٽ�άn#�XSj0;U��+z�`ۻ��rl���#��G���A�! �P`O�ۨ[@���lֳ6ح�8r[b C��x���u�xǽW�_J��a��AM�A�{%!��d�&T�DI��_��Q�Z,��l�Z�=k58pEX���bP�z���^dL�d�jAVa)BN�m1�kղ��2�ܠ=[���l�qƋ6�w� ��m�Z���h�Q2<���l���&!?.R_m��Q���z�w��BO�a�;�!�QN�a�I�����͔�:��T���?�S|�*gU��U,� ��
��	�}�OD�Qj�j�W��r����_�s�Zob(��f�'�=�`"��%_g�(�zs�b�Ծ�n�
���ڵy)��)>:Nw%�%�c�kOC��@�������S	Tt�e�t=ı7<O8��'&�*Ӄ]����{�����Njؤr�3u�_k��S��_M.�����-/ě)R&b�~��	Vġ��zn5`]�@�HKe��賔��y	�L����4\�
M@��H�h��*�����T���%l2vĶ3��[S�َ�n(K�`$c�I�
�`E�J�Y��s��N�Q��{X���;+�v�:
����,�� `�X������I2ER�%�V"ɼ/�+ֈ�4���э#al���!�iw��Xy"|�sw�iq@D	\���t�~�"��EЃ�7��g��(e^�}$�������O�u"����-�{W�)�>��1���mS���A��VH���*r�㨿!�Lm�(=K��ȷ�Q��%&��V�U+՗1���O���@��'�-F�m�Bh׾ۿ���'"λ�J�:�_��)w! ��"a7�5�}:_6����呑��my�,��V#�(���໻��l�XPY�G��N���SCe�)d����_��Ȓ6w�]���K(�ţd��᡿����81Y���}t�;�T��FH�|l	�
�@L_�L@��+��.�-^���Q���u5"��U��X开�f] Q��5�1iW/>�/���饀⋊J'n��fM�VH�W��c�U|~��+O�9B&��_�oX;��h�t{ף��[zWœ
C^�q�}/���Fg��|��{M�%�zU!_@=N�$��""2� �l��"U�e�wp-UO����r��S��9o˖���]©�|���3�H���]�m^��l�#���,����}>a��f8�@�N����.�LV����	b�S�0�.���W�"���e
$u?�ȓ2~�eź�$Vp�_cS�����qr���؎���g��եi��+�'�8�D�@ݏ�E�
<�zOI&P �tz����os%0ܮ�a�h��#S��#P1+���=,��َ���N���4&K���lJr�LX<�����R�s���tߖ�=��+'�:�%������C/�p��f�.�p�������8����������*O�_�;ه�Q*O�䴒<�b<���h�,��u/~���䐉G�B!���뙆�-c[�է�zg�;�H���uN!���m���zu���x]ۛ��,��;G/f���Rx{�嶢�lf��!HͿD�գ8qtjW��{P��6J��ME!���ȭk#�%�*g�_�Vsvc�q��ۉԈ��{�r�Ƒ�h��XV��y�s��
:�7�w𵵾	�<�ŇFC'��x�����+b�3�e���.7<ul���Rk�i�T���WJ�Ȥ�@2��r���/�#��.���Zk7�����G,��|-���(%�p�c	�1�>�`��ܘ$�2���`&J�Șc/��D�M�׉
�`jVۭE��`����J��v	��^7(��q]9kCw�ehr��y3j�A�O8(M�Q�V&!Ъ�j&�ځ#Ĝ!:��U�������FNV�������MB1�Q�[����_"!�Z�J[yG�}2g?;����î݊�J��mG\~
��BFF�ZK�oDzҾ1�7q�+�U����TM�7�Ma�
F;�7u3�����g�\�<L����dWi��Ϟg��+����,���R����"�N�2iʉL�j� ���gu���	֎��
�$����N*��b6_կ�֍�W@S�Zo|�d�Pػ�9"�'A��U�@	�����'ɡ]�Ms��F��w���OW��I|{�(g�^��_�_��~���e����"#A� ��E0�[.����]��"���� 19�X��p��K��G�b���Ύ6����������pUHSS �.o<h�p���q���2n��7�_����������7�)ʯ�([����v��MƢ�{�r.���$�}A��OVA��Y�5޷f]p�����O�U��vM^�9�z��|�e[`ON�tк�f�Oe�wT�I��t���Z��<��vǉL'${��'�͐=��s�of�I��Rq�6 .����p=��
@k�`>��D��������Sw�8 ��=W^��WQ������pm��"{,�[����H�ь;�#��[13!m\�з�5x||s�(_P�M�m[�0� �f�ٳZ�"f
|9�k��@,u+�ƫ�F%��S�U�����Dw�l��W6���}e�cU \�W�v�mU�k��&|�}��4E�k��V�c���$dmw����l�h�����ĩGށ���6�w�9L�������i�sDL��
hK�{��f쭍%���:�u���%YR_���KR��8�<�(j(-hhq��;O�e���Y��$:�r�V�o�Ng6�{�+�|���mv���f�uM㳘�n�b���W �eY�W�<A@b�����ކ,"���>���ҏ)��3)'�ҡ���D�s#t�0Xk�����]����M����f�Kz��Ќ�I���<��E�ck4��r@\�gE_|�m�<9g�A�Q�U�؛��ûE�#8V%ڒk�fc�ӂ%|A�vX]��ad]���R�@@#�,Ֆ_��$���ͬDu�sM��� �.�0/��m'��'5zkIgo�B��8���ĴYh������Mt]bCr�~°x�MQ��^�(�y�{تH��y1Hl���1܇Wuz��P��O$�����<���*�M���8`�mX�
n���#y��FR��v��0��� k�(�tI�{H��
h���Z�P���_!�d�'R�/
�tqV�Ǝ�`ip�1�ԉ/��-�/O����iC�C`�]�z�0�B�h֊�'d���;`�{f�b|D�d��I���GO��eX�����$j>�v[#�p\�31�Kr
���SP�\��-D�U�e�eʘl�v������<+�Z`?]�A��r�H���w�mf�&LZLʹ`̕˝�gy������2G��۶�Mf�3�}�"ថ�HH��"+y�	�v�a��32.)���7Kf� O~La���=+2�ɸ4��[����@q?Ei�.đ�ϳ;kͭ�%e�:���~���C�gi�βN����~�o� p�X7�	�� �a�i�4�5*�IU��~<eҼ���{��~6aO�Z��?'W���ۑ��mǔ�	�OtoR�H�p��T��m�y�PZN��<EY<g�*B�zB���5ISH ���+^�yD�ȑ�SU0���.��p-˗Xp)
ꞫBj�)b��Cʗ)�<䅔�����Y�#12�w-8���I Xӑ�F�#�M(�1�鹗Q0��l�n����[@V�cJ맦�Q=ىik�z�B���ۃ�hk��UZ�M��&�S�)I�i�A��>O.���'�Q5*��4�O�������ԧ�gڏdIS�������g��&��I�[��8�6)���x���-wQө�\��A��q)
<́=�ި���2b��Ś� }Vj�*M���0�j�q˩�:U��{@ͻd}�w!�u�eS�6�h�ЇPJS|��n>��� ,*�d|�B�hHU_J� ��'��{"3�I��j�h��w&�A���bM�mܛ���M�$��N�+m�n��Ȭ���j3Z�-L��Jr�K�\��ZނDu8_����1�Ɓ��F�i��]FML6�`�B���o�Y3j 9	q��W�R�}=/�&��.���{E�g�sn�#�ZoI�;@Ʌ���`c�TP`G��4Fx ���|��1�(߬�ޗ�6�?T&�c>��]<�1ɹ����L
٠d��J�Z�J&i��O%(ߟ����N�Һ�O�JT���-n�8H"�)�_TT���s=,��9��y�m~|��.ma,����+H�eM����vyr��M-�V�I�㵏#�ឞ��;<��M������<yf�r$���Pe%�d�Z�BM�N����3:�BQ�1E��]��-��,RM�G>Y�϶PjW+4i)9�;I�ULr��zyu�R�́9�2�����7�4���ͨ��ch�F�ԼB���㓓k�VR��Q`�m�#<��[Ǭ����Ԓ�&��A�1%���h�-�?8�678����9����{��v�9G�?�jβ���(�
�\���󀷫�dw�阵p�nbsY�jq�<��,�G$�*�?�\�Y���AY�w1�x�V��~�0����X8'��tBB�h��bA=��A�y���(iB����=��-deW#�����OPz�*>q��*�Q�zb!���E-ݕ�����s	B��&�+�Ua��4��kTӅ4}5L~� ���VaM����Dm�����Ξ��h��rR��)�H �s�J�t6&�=�h� ��WcNr�W�i��;��i|�8=aj���ԙ	u���ϔ�h� 3�_�&l���ؘІL�k�-6�Ծ��q�d��0Ӂ�`�7#�3��I����FZ]�]Le�Y@�B������<F�q+n�N��l�� G\߮|!�6�Q�:TM���)�P�M�% ��}LH��#԰�=�G�JY� �[�p��T%iEˢ�\R��ۭ�h	*Xy�7�ѷ�����ڽV�(�u��ɩv�12��4�n¯n���#���_���z�MOϱ$��)�u������ cq��G�����-��R˽���[�+�\Yʎ01a=Wq��vf�|��Mqu��� �TӚ��R鱹�K����3H#(�Byx��������Y�NQ�Kb��ER��8�d\��m��DEV	HQm)�U�5٩&�HqHU�"��D��=����2 ���Ա9�秼G-�k�_�,��&S1,����[�GQ8�jX�9�@�p=��	��k��EΡN��I�S���u9���9?���U`R-n�#]�t�*�� ඪ�O�<��Zfj�8���e�ZU��kڤ�[��oJ�-<�ɶW4<:5K�*ĐF8���e�XȈ�[m'�:%t6�m�*��	zii�`���P g��*5JW	�u��oSy@W��;��[�y��b�+�7�"zE�zԢ)U7CSm�Nm^��z�茾�O�R< �8VGi�)):�Q�wvx� ��Խ_��oGjV��V&�R�R��G`]�
B@9��f���y�����q�n=G��NɼXY8H>a��u�j��8	�������$�Q>i9 �<	X'�7��w�<�xa!o#��q��J��Z��\[8t�*"�+�$�ߟt
BPmm�ֿ�8�T:t�8=�>m�1�G�X������C��Rw]V�q'pM��H��|���IB���D-�uG�pP�қwzBk uQ7�%*�P�z�ő�.�R�/̐����WH�c������x�'
H9���@z�@YVm����$��q�hSjRT�6�_�qs{�A�R�nE�Dro�-�� �$����m�Ѿ��pH�+U�${#�U����-�X(^*l�B�#��4R��IR;�[��C<�+��sJHM���^����h6r ��X�+w;�	����T&��FLi$R.|`XK��d��|�ĭ��nVB��#l�I ^���$���J;o�E�[�[H��#��'h��z#�����j�Z��o&WdԩR )G����n�Q\�|M��h��ٗt!)�����6����I�tC�&���+����[")�"��P� h�� r�Й�fĆf���t)+��a�8�t�
�k��1 ���&��1ۄ��.%�Z{T��Tن�4����
���1��q���nC�7J���w`� י�t79�+�mT�����tO_���RW;4��S�*������)�����z����h|1�����%��W@Iu��'�L�\o���Dn;� ��M�C�]����-� CU� ��96�o�G%f:�=ÔH�i�J���Y�k+p�n=þ��CA=�jj�4I�R�ˎ`@9,��Y��D�9r��������M�{��� �:�-Ub�Cm�H��B%�F/pH�q�Z)�i�P�S��4�'�j�*@W�y�ߕ�-cH�ot�/	�����mgt=W��iM��eA˂�ɷ��ԚBz�*��1/5.W��ʯ��|j�v�E���y����x��wX��x�B�,4�����̴����[M�W�>w��X�L�6"��~��jZD�~N�%մ�OAQ<�X��GxM����d�ui�����E���×����v�B�Y]��*�R�L��@�g�<W�O��|H��ӵ��=7<f_TۋD�	R��6�R���[@uZ������3�w|�z'JЍ_7.��u-�-m�#�P���N���4�5^�R�2��ʓ��T�N+%`&׿X�f¼��b.�������8a�w�D�s��`��#׈ �Z�#�c���I<o��o�j��Pᕤ�  ��,':'�O[61��)Ϫ:*�@U%W�C�4̻Ȗ��%(�X;e۽��7'��G������H7.ˏ4��3��I�M�{���`r�����#3L�m��P�(en ��v�T��{�p6�/��y�v}��i�^N˩���-K'� aWJ�WQ���S����^ۢ�E#GP�4֡�麛s��{7�{rIQ)RE�!B�)P�Ův�Z=O�+R��NHV���[�oqn�ؠ��'��#�dvm�\�>�G�~��N�6E�N���7}n��U���{lO�%�Q*��cD�N���?T�s�:v�Cu�Sf; ��R�s����Ďp�����$���h�2���'L�� ��28��Bo�,�Ч諐6�� >���	���vc3�N�5)ڴ��'�<�m� �F��rI��Ď������e|���e$ �� 9�(G�I� �b!��%m���Rm{�� &���\\��&�II����%���O����!���s�q�z���K`+���Ģ����<ۧ��mt2bV��$��e^VJe�-��K(�"�G3�EkK79ʯ,� ����ڊ�@m�is��;����ߕ���$��m^9�5� �O�%���P�ȅ���@�� ��.�K�G|��A�*�vN��� �XOu~�i�O���9<J��>ZŇS.�a#�!.��q�(5R*L%-����HO�K�n��#R	HV���[���Ҹ��H����&�(k�LJ�l^\Bg�"l l<��ҴJ$�=/y=<)#j�y~����XZ��������iq^�}v�3T֛
[��A��?lW*\X�J�g�Ӄ�m���4uZ(;A� q%&�{D|�(�y�����\'��R�����p�������-�9��U����7O����7(�w�#�}�|�[u��B��]��ji� ��o�A��m�SU�4 3zk��LC�n"c��}ri�<l� $Ӕ��8J�5(�c?�>f���7&� B~��c��ԜA�h�]/W�ܫ�?4:���ۄg��x����R�͕$,=�ǌ��w�*���eo�_�4��ɮh�ͥ�\�-�E!���
��v��	� K�^?���<hֿ����?z
�5�sI�w�?~z<��|ԛU�
���V�Z�}���g:�BJL��u�}�HQ�8Jo�~�z@��l��H2i�G|��� :c����4�4��k��F�A�[��l���F��N�Y��J=��x�S�$���(|���{�NSV�G�	dj*rP�n��j��e�p���!d�
���� � H��k-]/���mҤ��m���c�a~gh7��W�NP�����E[&�?R��5-4����qI�e�4��\<bYMj�9�S�:�[��q�XAG8�p�7A#��5����_]�s����_߃޳�k�F���HsTɼ��AM-�-��`���2��K.� lJ).�����$8��������#�J����n�R~�D鵁��}�BV?Y��J'X��+�Od��ik����dj�7*�«b�
���m�8����46�V�X������qP����{�,��b��v Y�Tn֢���8wһn� ��>�?gU���'��x8 � � ��*�N�Ý2��� +�C���]�R8q�lq�b�0���D�q����Q��7'Q��..R�b��*�-��4�$�,0���� ��V \s6I��!j����6�?��zs�����#v����`�H����n�\&"��� ;�;�a�h^��.ɶE�NN���/�䇥��tZ�V-�$���u| ��Ywi��?eR��B�A ��55��FJ����N���Z2Z���D���Ęt�K����l����L
[8���4_�٢?ȩ{u�]_v:���yb?ُ݀#��M�+� ��*hX"��p�� 3�;��Ɇ�\(�V�}�!��}�����i�2�z\I	�֤4A�_	�bh�ͮ�,\\);�%��T����N�����O�"�Jo�� êe(�\�M��g*�6�g�y���|.�C�-"����թ��b��!:�Es�B�fU�2��'�V��>�R��e��M'�G��1`1�O{Z61�
=�ec�$�|p� �I"�1�C�D�_B�
S���(�qQVz���τp������{r$Z��R隅&F^�G~a�VCaH^р;�43|;S�+NNc�j~�T�zs���1!�������?�_)��GQ���Ui���)*]�}*6��(�9�j_y$�EJ�9χH��- �Q�؍�]Z��ϟ5��xA�~$k
~���vm>S;0��Y4�ir�֣�)�>�ü�ARUef�揔{�?�j��YSR�˶�?���*#��W����߲�dy���		�0뙙��$[�yd���&/�8���Ӓ����&6��Yl�Z&�v� �.R1�q�7d��,3�3]��9,ӛ��M�*��t�*#���#��%���/F���f���W�{fX)��8��Ap|c���u��\�)�2�IP��H� �GG��K�����g1�A��t�MI4��8�K�L�ڊ�E����P�TH�x���Jj�i4/غ�;*�<��)jMԥ��P
��Ty���P��2�!�-JHY�S����÷����̜(��6�XF���Vju��d۔�c$��C���+  N�z����6�6�l�̻M��Hi��%	�B�)_YW��S`c퇗l�gV��)�SG�"v�'�$����æL	� B�t�'�L�@m���Qdܐc�b�D��K��F��A0$��"��ǉ�ln<������w�$6c��d'�|.�(�du���9�@$$q�][��v�ZܡDܺz�<�R��E�
9�Bi6�� �@�� X�wB� �2 7�C���������@�:7��^�*�T	�ͳpG�}tL�@qh!l\��ddZ��* r�8�G���)�zBkf�ߕd=<ͺ�qbNL�85ɂ��<a�ċkE��p9ı�"�&�v��q��	�/
�5"S��!��	X�2b��i(* [�#�d\t=��G��]��@�NS��`s��)6���:�c��$e�9#�: K'��y � �@*Y$���dzO ��@��N������}�S	ܠW(��� �O�Nm�D���ap�M�E�(�`CLnK�pU�ʦ�I�	����z�J�*�/8�)0698NT"eոX���V��bpȔ���{^
�=�G���E.��rû/��[w(��}ug�%�*

��#��]7?X�|TIK���ό
C�6�oLKd�#��;�|�o�Bo|TZ|��\�c�L�>�����O%0�r@�Vo���g�Ș_�;����zϔ$�L���$D�@6N!v�F�I���W$�2C�cR�� �0幉�Za����äJ�2}�e�[`{bP�\������o+���_]���o�C��0�ln8#�6͈8�J#+�4��B�P����r�ڐ����x<��-� ��  �$h�Dd���"r�I_9b?��ǾL�A%?�3�6�_� �2,rRE�*E�?�,���B�Bw����0s;R���� ���B���m���{ĭ&:I<ф�Ov*3�ܿW�9ǧ33s/���@��0 �I77������>(�ŽPl�����H�cr��a�������dM��x�!�*9�	�m�*���$$r� m��������:��#$Xr��)�EsҪR-�'�y�d�{�mE	�[�1dѺ�Y��	�Q�����H��Z���U�v���[����JIޒB�[�9Y*|�Eu9J]>Zy�wL�,��I�w{���ɀh_[�j��x�VY)����[jTl#�Ch骛����b�C��Mԍ��t�v��OM��6P,�{��eԭ��*�v��K�Q���>�HiE@�7�+�/�;\��HQ���Wh���Ed�.	�@"����x�����}Bu3�zb�����ЦB�yJI�����N�ə*E>Z�.Hܖb�rܣ�+�LI$䶂��ڸv�mIS$��d�*�&�P�<ԫt����B������tr/:�ϒY\����PK   |aSU��|�`  �c  /   images/290656fc-115e-450b-8d33-ab580af06883.jpg��P\��.:���0@��܂3.�>��wܝ�AB�0H���>������=����[�^�[]���^�W�ղ���0��
 R�W�``` �&����7J22�Z��J���
 �G����� ppts�R�~��o��dnu���W���?8 0��i�?�3K+�����ovs���_��1��?��?����`W-��8�/~c���`O7g�����-�]���b1{w��7 ��������� (@� ���`����=�N ��% ���� @s @9��:��6~ �F��]���������G � �� H~ 8��g�������e���o�����( ο���<, d X��?���˰���`�=��K������	�?'&$&&!R��R�S2PR����ӓP�dzI���������b?�&x���������5=t��b�b�cb�<"��$�x����$l��f�G������g�rD LL�G�XO?�~��������sn)l͗<�.���Jk%�1�~��@��/�
cֶN�;9�)X���
����寈�����P��ď0��K���6'qy��a��c$W/_�|����譏��(ڜ��T_R����x��.P�`�\PHU^+�n�y�@<j~,�h
�p'#�fkf�Z��G��sj�+�x������1����>O���z{�����IS2<�6_�I��&$���a݈���D7�����x�e(�Fx�^�P�Z�rS�d���X$�SC�Zdl'�K��Z>o,��d�R��~��<�cA"�B�"�"�o���m���Aa������ы�t"e��E*�zy_`_�z w��A�,��������jAxP9R0%�uB�'F�d]Y��.���Q��}�i�#�rDډ��s��t1��#��*@�(c�_yA8f^�Tj��qK.��A����ʛppC+�_��>4i�����m��Ⓙ #�7�Y<L�A�^�7w+K�|��d�Qk(ʁy���n��de����|*e���	R��8��+n���pq"$R܃���|TW����~�?�Q�e���)3z�F��Ŧ�`�p�i���I���p~Ӟ?r'uǨ��ev�>�yi��֍ţĄ����tQ�-¼n�|>����׍s�%dM�Z3����.�0?��)�ۃL�8�ZU�hc���`������ �֞$�[}�)�V�&��������w�]q���11a�쾄�qr������e��1g�C�ۗl*�s*MǊ��3��u�H��S�:V�-aK��{�_f���D3�rVNm���`O�x�;������/�B�����0?}�y��gb�$�"�6��z�:̅�(�߱�%�2�Z����#J�}�p7�&�X�Z�P�%��uڔ��)���B��K����(/c�B	�aٱ����Np��$��=��]�4�ؙ�O�U��t1?�"E_FDSQ2(�%`MÚ�G�*�CJ�}�c����3R-����Ue�/�}�X��2#�R�++���A|",�9���b����^p��<�a�h�N;a]H��ℯ��-Ƞ���.�-��M;-t9�<qH��#��9Ϻ���{����(/-�Z��()�9t��,kޛe��{��6�����X��j�R��d�9���p*y�]�K#-j��b�N-#
s�4��S&H�S���!�G������sƍ�Y���)HkԳU.۴�%�ɦ��U���������1yq�e� Z�62gu$$��0�y��Ў���l�ݭ2���O�t�!����~ki@3�R��|��s �Q =)�
[�R�������t*ux0{͎zA��?[[[LXzB��d���S���.��OVOt9lF�Jx�]��*�~����UIկh���;�u�w,ٖ�0����E��w�9��`V� "��ͥ!���ڱ�ƅ�A�S�e�ں.�;��Tˈ	�qT�j��aWq�	M�櫐qoc�%�<N`;�ǿ�#�/�9e�j���ҰA���*���&
ӝ��$K˛�f0=��QV ��8E�Xd��5!�U�+�0����iʈf����H	��먶��k��5+�Z1�OF����UG�56�Y`&���\\��M!Q=�U&/�񓂿��⟐�R���1�f�uY�6-�q\g/��S�f���=os��Ӓ`���002*}��>k>�x+��ɤ7�-��lӛ�����`nwE0�CE���t<���U-���5#��H*#�:IA�lrw���I^7�VT�螪��Y��;�:��S��ڑ}��+w�܌�\�D�ß�K�=�c�˘��+�9z��VĲ��Z�4Vq�0k����}��X�����3�$ w:���S�|�$�U�p�c*-�Yk�@cj�d�1C�Ůg��}s*w�y����\�%`ܵ���*UHmsl���} �TF_Cb�����?��"h�g�f�ț\w�I��Ŋ$ȉ���g��g�Ua�:�'Mu�Fq��aD�W�[�=��0�ZVT���o�~�^�j����s9�Wo=<�\�J�z�yLKJ�����fz�%Lz�~����}���J%�+Np@E��ɍn����"�v�J��<˛��D�IΒ�Qd��^�ǜo�PV�KJ���R���uhpِSk�bv��9s��A�u��&��A9<Ԇ�q��n%:5m:?��z�EL��7H���WfXY���B�!�}�92����� ��>��9ͦ���I侩�����T�j���3��2a�4��K�}�0|1k�ܧ���Z�V�H�;�>��W��J{ H,߯u �pq���0{(6��"���+8��;ν�kC�;�D���c�Ю]Q��m?#��^��P��9�E�,���ˑ�Q���o��(Gld��ɹYD�̺C3c������#�a���o\F[�)ڶ������r����n�D���@՝�e��o��ώ/I��2P40�0nxS�����UD~�.nŉz9�w�=�8�>�uOk��Z\��?d&��3\BТ.�=��"*o��K�Q���E��6n��T"��MG���O
��[����ӓ}�����)E�V����6���2�Ȝ"���Ūe��'�.� ��=g.��"�p"zFVs�� ��TPl�p̵��F�*��r)��c�a4�h��]�	�+�_?M���U�Ѥ��A����G����"�ᎁrό�ؼ��XY�6{�uAZw̯s�p��5��%x�JB�ᅰ��L�d}�QWPQ,�8n�w�aTAz�<�N�K|�RG\�V��(�G�p�J�Y�zJ��CQ�N~��G�1Uij���fc)�{~��
j��`;�ΰ�ӷ��rW׽��\��m��jƻq�'��'��U����,��{��<3�B~���C�7 �ƹ&�t4z�N�'����r���̦E�g%�r���$�~U��{ëE��h�� kZq~�;�J�[��vUN�ym������Uz�]��_�1UR�y�^d���cJ�ҧAW����U�2e?�յ�<
�sն���s�ś5��K�KS&���Si��
���v8��o���fl�1�Zt�y�mv�T�����K�K�B1����j�g�)J��Wy��k�D�D��j9�����N͌6w��v�� V�+�}�j�2t��!W�lB���Zb_�<�`J��M%� .}|k2����J�ps41*,����t�'6�j³�p� � 7�ֻ�XQ�;z���?�э�:Ao��5�DXоd����9�Q\{�'�mՇ�O�
ֺ��_޾�<�^�0,g���&>a�y<,��<��O�쫈��~��7�,y�����{�t5ՙ��ܸ��ۏ��Lx D,H�4M��`����%��Ɗ"~��g���#H�H��lU,��k��aώA!�F2YX#{�P�6D[.�y߱�9��D�ѥ�-��a�J�X ,k)�)���>��T���I��T��Px6��L@/�g��-k��吐��'�㭵5��S �����E�3���Н�V�(���Q�(YY�0�}��#�r*��=������������ 	���"{��p�y���n��c�f�-��g㙮լ�
�ˎFnE�-g5�����b�zF�G#^r�lZ��s���  udc���E��&k��:)���.���P����OGǷ�UEO���Qhr���hJ�_y2#n-�������S\:<s0�u)��R�h�ڪG+U�2/�K�����������4��xzO��e�e}ٙx��9�;�)v8jU���<��Z�1-+��$���Sz�ɥ��\�ķ�I�ߚ�LC%�Rk`��[g�M��%���ZwC�
_��l>��Q�۷��\���ߙ�W66[��9} �m�V������KFU���o�um�\f���nܠ���"���2n�������HģH�Ӻг������ncYIY�nkb�ڌ�X������k%`�=��������5h����o����#�}Y�D3���Ε�FO*N���g�)�M�P���4Eȅ�TT��!���V�۱,��~-��WY�W�Jr�Ӓ��k�)E��8KNP U~v��&��#rD:&�T���V~%��tq�q�g &�(��b�s�v��r*�~�$x�a׶���}x&m<C{B(�p��\8&�ե��A�<ެ�d�F���N�ņ��&}�1s`}N� �;��������V�w� �8��
 �j4(�MC���������I1�Gȷ½}>��&��������vtl�T>���>������F�d�ء
�(YH�����`���%d�f�+
����k�t��&ǣ���!&��?|��<����f�83!�߹�0Z}m,_��F�}���7�4�.,tة�����C"�E��?uk����^;�#�M*3�Y_z�M;�{��	����'��*�]�ԧHfKH�N�)��>r=9���ʕ�:��
6�P]��%�8��3�(�a��L<�R��v�aGHa�9e�~��N꘰����|��u����u�Y	��������e2��8I ����01�Οy9n���?O�l�c�g�u�ب���{����y�*ig��
��:G�9���/PqE�;o���\�(�6�P*0d�,��XWs�b�Zl��dK��\�,�N=6��d�Um.����/�&Q��tǴy?l���X��92F�Ϩ\Tey�fEn��@	������͡�ӄ�/�I�Lz�����C $SW�{+��Z���Ӏ�j�D%��P"���.������� ��w�l�UIKU�'���n��J�����l��N0�	ie�!�׏"\v�5":|*J�0Z\� �_읻������W��/ih��ي�6C��9Q~7�J���M���c$J��u7��e�_}��?���	_�l勱�<�֯���El��k��?ͳ�t�`.���A��V2�~�O�|�xXnD�[�d�����wg��_+��'Т�ĲL4��AY9��W���%�HM��ts����&���cca�J%өGl2�@�,�������|X�3��YS���VsX�zm2N���	�I(EЅ������~L�׳7h%&��g�Z"��e�!��d�T���S�|��Y_7�~�Ɋ_��k�i!���P�Y��z�:�C�6ź݄��B�}U��������}���Q�pU�\�8$��^�H�-;�c;��SP~ۍ��P�}B}e/�5�z�bBYr��p'|��9���|��F�?~֝ؒM:��f����OiL��������,3�xxO�R:�f�rF����7Jz�����{��M�!��]�K�K5}�����:��W|QM��R�ǖ��`�V���'�.\^�����Ԥ�=6iC G�'~���\
�JN|��K}jQi7���T/
x�[�=Vs�a@h�����9��n[��h�n�lT�5K��uh�Z�ѡ�n%�os��П!�99�s����K\&A)�¦��-;׃1:��F�=�c�Z5*�=�&�Ф��Qȝ���@�oM���JX�t�6ю����>��ZN���R�3�]���/�ϭ�b���U��V`�����µvI��>Mbr���
ʣ�n�WKYf�ӑ�49��
�����o�#�F�b�u�3�w�i_'��T�6�@[]���ۑ�ϡ����Yŕ���N���.�م��w���Q�2kq�	�PM�h�aO�5N��ίs�⮣�DI�,����F*8�l�'J=42�t�{�PZ7.�pF�L͛�ݏ���|sN�@*rsZ���,K�������<I�k���f'�7o�m��r6B�>�=�T�`�y��_����a]�S�|�Q�қ�ꆛ��Q�<z$C���e�/��6��ė�.�ђ��4D�V��[�"��u�I�̟�$d�Qw��5���(��&õ�o��V[K;��?�)�c�Ħ�{��	�qT?���~��[��~�1AF&����x�G�X�"�����Ljm�}�s�{��4쒂�,k�:m �Sw�~��8G�T^/��HE[�.;��?��D���W<�_&w�z�a}]��@���͎��J�0G���`2���9��ˉ�K�����-;���!�*�*a�j�2!��O��z.�t|�lO*�@9��{��;8��
'����w^3�A��4ﳽ/��*���	AЫE�9��g6�^�ﳢY��_�����~h�\3BQw�I�Rr��&_��)���7nڨ�g���[Sr&��!E��^-L�O�Q\�����j� �U���7͗�{ث>�d��"�v��ʂy�^x�c��ף~�!<uO��qu��M3j�g}]�7��o�[C�v,oЖP��-y��C�I?rl)��j��p$���6׋���4gM�֦������(���)3���2AME�f1��[�����e�VZ֎�@�j^>)�<.��:AI��˗t6�C�`�Rw^����=�I#o���-zC�*f�B�����|~����`I����,�f�n[X�-�5d���:>����f��`��Y�nעf�[hf�򸺯i�$aNA�1���Ơ	ݧ�Yfq-C������M�����H����T�?F�Ǣ��?X�ӱ������������.�K�� ؽ˟W��������nmB]�ŝ1�\<�?ׅ�F�fg�;+TCZu?�D�G ��ijgX�jd�[ޣ�j����@��Q/H��n���O�⁀�wn��<��/����ݕ��F H�g��^�QT��dB�/x��z�H����Q����v�`j܁Z�ۺv��Q7��x
�?�S�	p��K�%_���e��e@+j�t��?%�"���хc��;}� �b�,哷9^�q��;C��د�8�[T�W��D�|��oJR���na���GD?{���w�?�V�w{����< ��Q%�W��!^�	�1hq>m�:��-hIpAD4����:rR�wp�/�p/H���<�Q��\$��9	���ǥ�꛲<-���e��ؖ��Pb>ÚG������B���X����/�����Ws]��stBǬ�L��n�ԡ��aIS��0l�o֝6�o⟨��C(��|*V61D��0�m0Y�E��7.a�������&��e�|��U�x#��:u�L�^�dL��M�ִ��?���2ݤ+�Ƌ�)w|�5�m7(e?JK�aΞ|���J�=��Mh���PX�Ӧ�-E�-5� Ȩ��"�k<��������?\\8�A����iO�~<!�0��e}�v�O �o,�uCX�3�+� nCC�rմT�eW��[ť������J
��K�lg��O/�9T����!cƈ���~-�vK]+!�v���EC~tk�"0���t+SB�̇��~��}�H��O)L}q���^�[ ��XZתa���D�,�4��6��%:\2TCy6�^%Yn\y���HTS���tU�v�(םc4\�ز�8�.��Qb�lx6L�|��l��̺�ʚ�4��6�͘�V#^B< �֚<��ٕd��CLb��e����%��~X�C��S��F�ɕ��$1(�NwA+��~s&sS��%��G����6V'��:�Ԇ��AС�r�f���J��U i�T�H
/�Nﱟ/<��lW2L��e�e�uGW�l~pu��W^��K��omK*�f�)��d}�-Qm^�*�iZ�;�n�+z�. �~M?M?s�}�Ϫ���~����,@o��dQ���~V����+����K�o݉K��z-��P(��o�r�tb"/��D����b���iQSU�[��Ԝ�m����;[��SCetф�N�R*��F�^�H��R�����]�\�4�8CZ8ZG����3�voo���/&��hO�t�`���@=L���o�=��u�=b�i�Tu�,]}N���K1Z��D_�ϙ_:ps��a��?�KR��`v��;̟�d�|>]s�6�r�Q1v[A�q:OJdl<VM�\�����*�=erHh�	b�$�:�~�rH�_����b%1a��M�@*�/&����ַ�,k�W�z;�:=!O��գ�������)���*2���N���-렒���ONK��!�+>T��j7����e�A�a�2]��?ȈŶb	�[�A��|ב�=Z�%�S�����.�G{�����y���1G/��9����������$�tC�U�7d��e�E+��e���X��ru���Qܿ��
�[��	>E7�_��M���	}���Ǯ=����5�?V�neIA�S��(��9�B�~:Z;/�v~��)�k�0���� }�b��������Zf��), �s~�J����I���́�� �!>�Ϭ��%�[�:sI��ykm<�Qat�b��B�O-4R`Bv�ʠ>ݔ����D���)
5�~�['^��P{�	3oa`�%�\KW7�A��C�
NB,l���O)zi`G�����v7/Z!�38�z4��6S�կJ~�aDr�V������s��ܑ�ƶ��ߡ���q����)U�rr�h�*	�sA��K�U�:o�l�|�5�N�)�uQ�%�r9X�!����q*�u�����`���
ip�Tg�$`w-G����'D>��U۞j�e\ܧ;����;�#���P�:���W�CoǔWm6�IP���_��gzǄ34�χK��7T���Ф�Ʈ���˩{���ϙ�|$��ޒ����m�)�
n�0~߇�my���H��*�Ǒ���C��> �zB���X@xd=��,e˳�T���<�5�KE�q��YT�1�� Ld�ux���d���v���45=�0���x~"C;�$��U��RR�C<�=�Zу�|�v�'�u9��`��{��f�L֥.�)qF�K�u��e�����[k�&R�ۅ��$缔qr��f��wp�h�uj���y&�L�s��_���;g��a�wQF'ݝl�-Ϭ�0�1Ս��qӮ+�+)��'����c!N �����[:�=���K���U8�ϔj� L*�&�0���Y����I�m S�{�y�5�w:�A�����<�+n�)��x��a�W`�^��oI,���`r��U��Ekelz��[��]ś��m�
E��߷�ww֡�H�jb�4
9h�{*<���q`F9/����i@n�߶�8�� �SBs��< ��)s��|� W�eF�ui�v}�Y��V����bE��]�R?].��g�^�7�+��{RWEz!�e��XЊ�_�T8����[�t�����R.k!c���r_&�k^�����es�-Ge������E�N�%.���ੰۣ�ٲoN��t��}b�����-�����	�]$JY�~��.<�7���t��l5���;P���Q�TH��٪Z���Xk/q"<�^�(r2�d_����L(��Ht���ngy�[�[�8��� ֡Y�GM�EN���@���h���+!�ɗ��)5�R��[���0�~Y�����u�p2��&�� L/�/H��ˀ���� \�=K�����>�@T�*�,����$(��0}=s/��t3��%)���V���r9@�@���1��*k#���~(�*g�ꈵ>�@���(���UɟN�4���.��((���#�n�'����(fk̦���6��N��'+�z�����9��6��ͯ�I%�5VMHg����u��c!��W�o�M��hYi����:ds��S&i��+�'�k#�ن������1W�ޖ����l5Q��s��j8K�Y;�zc�w< �3e~,��'�#3�9���:��>���SS�����^�9Y�m:�������S���ૐa+���_(�bߐn�7��N�t�)ǉc"B�,{�׺�������Ȃ���q�{
ܽ���)�O����O���琰�@���
�jxd��Aq�I�m;!|���ݤ�o��N�r:K��� h0�:�]��L��2ss�$�?!����f�:V����wN�Bl?:7�|���8��]��n}�ky����,�ŏ����1A��L��n7
&��/�+I]QLք��ȃ��ߠ�ݧILoE��Ճ��z�M0���ur���8d��9��M�z���)���qt ���wǆy���i�2�ª����U�\�ylw�8�I�@��B�_"�O߻cz��i�aq�Ï��I��U��6�r&Hh��R�'~���T`4�C�Y�^�
���a��!	,����>QN�N�����.�L��r�M���u{«���$,�I�Y�I�΀�Wuq��F��p�%�GSV���R�|k�-Y�훭�X��VD��+�{xSD"�g ���&=:#�)�'.1��:g�I�����<Vf�7a^0P�����^w`�考^�s�Ȏ��0Q�ѧ��cN)v��!��k��j#h�p#j/�[�cY���c�V���%���D� ��d?��!�L;�\��R��>��ƾHU}S�\�EE���{S��,7q���}�L�QV��-s���������"��]�4�g�2�B��(s�A4R:��ߗ�g�]E��K���DM>�aG�$����gю��*_��h�L
���Ql�@������ᜅ�<b'g�YVQ���f\�K���m�o�~��
]�<9��K 3{�V��jc�*���:U��nm�������O+�d�����/�͸ Ɍة�}���XPO��+=���:e���6����A�Y�b���9͝s��Ա,.�..o7 c��xô�)vC֨ ;�O�<d�I����'��z`;F�A���\+��C�����uN_%&8��ZdV�%��	y��[�q���e��]��=��`�<8u�nr���uR��
Զ��{�����	T��=�9ý�A�-3����QX�����B�Xq��hF��B���i	�!��X)a�$o\��6i��ENY��}P��'��pϳ������k�"���H���Û5���-���"�ˬü��1˾Ϗv�am�a���=�ӭS|5);�������w����l|��}kQL�wV��1JL"�9�.�ϽA<|[���o���T��4�8�;���n@��wy'~r:]EV5p�kˣ�� zx���K�M{9d��=qX�8������Ƿ`�k�`2�
~-<TW�3���˺C�M��G���I͘�c�̐>î{6B�x{�������祱5��*��YQ���l��z[��e��^����4�	ż>��]��������ۓ���F3ᘡ� �[��p��J��fB�~��@���ݕM'?����߷Њ�e��-=�($m����/2�>��c���&Q���
7�j��55	9���û�X
��k�f�!ض^B�e2�+��*����8���Y_x�=�f�%�� ,�}���m�{[�B��'�o�o�
d��yi��{:5�Ӥ�nf�B���I�!i�Z���>�[��h��F�y u�)���<M�M�� ~��d������},����$w�"�<��3>�S���ܟ�'`�i�"sWV�TV��t5�}�a�;�~ɚ��Pk� ���1�.�w�Yb�H�	|�ĉ����*J\�X��"�g�^*$բ)��lǩq��$�*%G�~Z�)0ލ-5�@+�;�u*c8eY�SY:�� 5qǁ�����2Pd*�N���ڈ~���Q�]w�Ƈ@��kf�Y���I��ă�&�^J gV����Q8ڝ�j��Ӣ�4y8:�_�l��1u�t;���j�QeT���65�2e�S��*;��6i� w�|pR���EEO�,6C�;(���52�q[(kU�l�s����`iC	�1~�a���'��ua�oI��^;|A����q6�����T�\�����YCSPu��Q��d����$���v�0����e� 8��q= r�y�f�
m����������[�������ׅ����0���?��}�R�pc���.�U�Ե�"u��)�����]&W#m����.�F:,�%>���Wܧ�TH��jmŎ.d�v�iwE�(ѿ���ʤYJ�6׵�r�{{��c�Hq?1�~��� ER=NYΞ��lV��pnE4۪Y�j��!\��)����R������@g]�����|������m�z�3���N�07����rv�jM�9֐Q2F�u��~]l��? �?�-*�:�'�����o8�:����8����N��aS��cV<�(\OY���*��$2rIz �����$�9�̑	(�3S�_�F�NA��ע�V���.;N+�&w�o�T��N� JF_�!R����AA�.B6Q���K���m]��M�m��n(���D�^:b�9�~l����s�	�\�Rc��ww�%�� '3a^ �ٷ��s�H,��%$c��)i�;�\�a62��0������
͍���pRk�>�h�&\;�Ol���m�o+�7�6498�	�Ub�T^���6#��Kn��Nh�Ăc�0�s�,}���^��,�eWM===c�'���1�����w�.2#� I!U�A�[�.u-���l�W���-un��S��% �lz%e�))v�|�Ox�g���A�I�ۇ.6L>dC���S��R�͈oÏ���Ф���U�T�DLlUKLD�mX�� ����k���WrG�M�C�Y�"�1,Y�e�uC���w;t_��Ϡ�Ŕ+�<���m~�_�l�)mX{���uB��a�}���$B��k��TN�žWޣ�D5�����Z�q�i��� �
r�Gb�.�('�P47��˄ۭ���D�g���l�������B�=|Fα��_L*����;l$=z x��r? p��>E;'�@	�Q�����ۡ�a��d��冷b��T�&E��w`��>��� ���'L�?��! |�8��8�ÌY�a?v�J�����nu{8K���M�����p�.FD,���r�E��?����U�#�<9<���� �g8�>Q{ }���w"�ڄs�_�n�^��""d����>�U�S��H6�sMk%��Ry����,.}-��$ٍ�(�����nޚ��G)DoV��W6��s׍̖Ҧ�4���2B!�3T�q���-:�hO��3pLI<Y��|�O��c�j;Õ�L�-�5)�9��e,^��/<Qo'X������x!��-�k��F,^j0Ғ�����1o�/���M�����x���F /�C~��q�U�d����"��8(�����!��	�\�g��)�	W�KPw��V�b_���}
�Ԃ��p�~�QRznx�SSLyժ/X�,���Bn�id$�j֧l��L����Uq�´�"��Y��Auv�u��+Pd=O�|@[�I瞜UB?G��e���0�Ud*F66�a*euc=�~�ͷ���{y�8>1�O�-�2�jn�V��Ç���T�u��L�I�u����r��������y��@��N�J�V��Ƭ��+؝��O���1���䔏ÂebʫEs�ÆKc�A�$�W砬�֦��7��ڒĥ�t��3X�N�h���̂u������j�v�"���պ�~:D��Rx�2#�^W.�0�	�fC�|�7��z���>σ&DM0�]�Woh��{�Jm��=�$4c���6k`�Q81�b�?�?���̆Kq ��J��Gm%:��;ҳ�\<��z¾y�5%iFX,���?���|����������HϿ[)/�3&��+V��H���$���M���]L�_�3�M��:�3����F�֏�2%�ۈ�)^�-2A+�A4}���q:h<5�� ^��M�Idb�`��5�Rp��1|:�vt��j[.3�q�C�j��[<�Sx��acQZjI����S��α��ֽ�3Ʌ��[z��'���Ú	E�®�{^�Gq��Ո��G���b��o��o@�&�ι���1�����2s�<���dt�b��("[z:�P�O1��P����m��TT�@_�������4�ǡ7�};�f�j,�d>��J|@@�`��ݫ�����4�Û�+oN% �|z���7�Oj1�s��zx`�7�ԁ���3��i���ٷ���JϘ|=R>5�e��^+�K;�[&�؁� ��h�sl8�K��d|��7k?;� ;�8��������T�˲/��ȃ��\U�-=�4�`D�./yj��7'kdTUɾ��~����~7zmt�7ý�V%Z5���+O���Ɲ�v�{&�^`���j���RDW�!(��H�f��������S�H[�����Ϥ6�Mr��`�.f��r�bu�/j�'/��ʫ�69 O��$k����(����ġ�]Fƾ�_LiR�w�&`�\��V��QG�Fl�Hf����W��e���z)(�U���Qf;�GHu�seB�rw�[,'���7��k���!���sWQ���2i�K&Jg��3F�w�]��1�.����¼�������EW��ޙ�bb�����)���z�-�\1���WhZ�x��a�������1l��e�n��*���/�gq��Py�����^�����Wx���ϻ���腲*wDɹH��Y~��;6������P�̩D�0e�UdB�,�1�������e���/�(�ѣ���ƍ~0��T*
w�.-��j e�$ˮ�n�i��s�ؙ�u՜��C���Yg�:y�=!=b����1,a|�0�Q�fH}��������ɺg��)fJ�B����Ѫ���cb1<�-_p���f%��� ��u)Q��B�xK����d	�A��M��my�PJv@i��fBm�_݅��O������:�#_h��ޝ���v��cgT��'
ҭ�Pe�Y���?��@+��㵯����0��o�����I1"�*���Վ����2����y"6��*P�g�焂�;D�F�Mׯ5�I_�c3_�@����Йt��P�5n�]\"]��,AV.U�ohD�߻g��3���9�
r�)�>�ǀ���m��3b�A��q�9��θ�p���:�=!ڔ�Pʔo���}ǻ��z:��� ���vӶΡB4Ā�&( �u��"�
� І���9�\�vm�U&? @�G�c�*֚ '�@h ��ѵ#G��] $��Om.zh�/a�|<	���[�:����e����CSlJ����.o�v6�<AU�wOX[�q�OqS}�rA�%�t uO3.J"�F�K�yIPĀŞ�`���˝��Z}��>ܠq�h�&FniTa���	�f=���x��D ��H
0k�!����>ܝ|�3��,؃0�b(���61�Ӫ�$X��Y�H
�Z���/j�����=��U��d�8Z�9=A7���{�-���sy����z 4��N ���-rof]�ZW@e��_�b�l�69����m�	"+�}$-���Z�wB���st#�uk��:!O�����(�}��>�&p�
��6�.�
"�鸅�������EK��{�����(��E���ϔ�6Pt�+Gaa�q�BW���S)�:�j�QV^bȔ�"o7 Thj�A�(�L��d�<�p	�F^�mr7|�Z�FdAaQ�3E~Oj��ּ}F�R)o��LG�g���U�㑈��J�5��T�vيom�Wν	�ڮ��6�y�Au?�~ $=����K1�����Uv(>�}��#�Pv���=��6�����^�r��� �?*�F�a����2dh�x����Pge#�8��
%	k��ђq�& +�l�&�7�]csw)�r���p�������E��mL�y�ȸ]+N�0K�|�\�����D��:��Xs/ w�k,�8�W�ѺC�y�y����x��a�'`Q�����~.}�mQ�y������s����آ����wF��}k�B�$ZD�0���5�E��2э&He�D�0m3A�]����%�ޢ�����׻�������ᬵ�������:;�e�L+6<&�c����5�'"������J0��X�izkc����X�� ��Y�����}��������{s��7�4E�1�U|�cV6��g�c(m�����T����@xE��0J.�Z�52��L�<)�ntZ4����� h�=$��f�j����I��P(��篫-Q'E��e��f��@޹BE�j���>w;s����s���-��o\���Z8���e84&�>*�l(��-���ɔ����Mx�(����޿�WR��ʂ�=>��Um�Yv������E�D.��Z���[�!r���1LG������,��b��Gp�O�G�1�y��b�����YQ�d����E�T���uL�m�g���s�:�\]��?��-X��o��)��n@ᅯq6�C�N���A))���<ְ폞23�kn�\m<�0!ΘA$��+�L|	����Z?��hnھ��H���02�O����mIZTo���9�e��=엯=]�鏤a� ����:�� �m{u͗�k,)-;�g�z77�Ǿ����
c��	��8b򡀫�6loM��-���{+ʱ����T����G��0T�>���V��4&�Id��s�ƒ24��x�Y�1č*�,+Tfp"���'%��߫ӣ,�:�{⬙�
�x�6�s�bfL������索�s�v�o�ڝ(�u�c�;�'��J���H�+x�6���ň����Pr������\7����q?�*�S�XH�,��H���Kx����
�3;Ӟ �3�U=��|�#��^FN<	�+�P�Z@Ex��/�;�,]g�\vh������iЂ�&�g?qI2z��=��h�gfQ�,w��ے$�XKm2-/�
0��F?�+:��=���x���y��/��+�-cq#�7ќxɈ�w����C�L�E)Ǖt�K5+�J��x�yzCT�v�1�@ןUj�}�d_��2���1����=�i�r��G��&�0�\��knޟRUo�n�:�tV�R.�\ үDV���Ŏ8�,�Ї2�&��Y0j��`[n¬q0�=�I,n-.������I�h�ȸ��\��\�H���X��uI��`��auQ�Oa���{�G��	��-�<B�I ������=5�nn��Sڠ��<��-O��]<e�uRJ���y{]�(S��2��҈%�<A�(>"ùI��ۯ���z����ݡU�#���H7}�i���Uk��񖆸@�?��d$�άa�Q5�����T�9�Zo=�n|��F�����8��~�s�@�;ehץY���MM��&�*1���F�h/0�JF�o	�Xo�W�Mt�E/� ����z���QiI<+~p&���a�xj�מ�:�K�X��+��&?�Z�0,Ӷ�v��_� ��}��N���'�CjulU+�/ж_@��X�W�ؗ��޲�@���\��0XC��i{�~�j8ؑ�O+FjB�{���z<sFEz�19k|F�A�;.�5�t��5e���vS��ؓ�ߠ��I\I�T��`�V�̲ٸ�Ws��g�u��OGiko�MO\��� ��4>�)�l��êf�t~
�R��i"�q���bӧ���%�:�l��^�s�쎢S+��߱�E��>�PeI�o�&���Ņ5s�:O~����^U/Uo%d�k�=`����dq�t�oɧ>A�9����{�:;�a<���	^U�TM^���ay� �~�/��Zn��E� ͌x��:R� ~�0�j��C3��p�[(+L7�nq�?�vw�� �cy�mƪ�!�Y��Z�s0�qi�~;0L��,��T�H���=��i��NQ
�.F���JIZ��
��e~`f/c��0����;Z	i�/��8��&��(�g����DZ[
��3뺅}[';;�L9�l7(f��)�GM�:��]7x=Tǿ�i�0t�̧f���֫���D.c'C ���@���۷���{�K�^�WW���d���"R�9�ɝ�Y�2�o"p���]^����8��G�d��{�ސ��F��ܲ�'3�v�.{<r~�D�y��)/�'�7ɩ<}��z���+�d�I�(��Pfl.gG�0���������UG�����\ ��&��U���:�[Y&��-���zh���R�G� ����$4��&�X�e^+�Y������ncɷqݛR�!�f��mJ=�~
n>��W.iGd��^U:��)��OT��H����m��!�M�o��T�Y;��b�v��.�^ ~��i�+���l��Ō��2Lg��U�۪�7��5#���&O�)��X����(WW��*���q��D/�[R�a��ξ���^�i��b^l�e߇k2'�j�JtH���� [MB�/fz�Vq&�O���g��W�����#�$/�I�U����+��Go�/�y��*��B����d��",d��v/���0x�}����~���}�W5))���wY~�7i|�Ƶ�~[��ҽl�����& ���<��w�_\  �OTP�z��,�Y`��2��ưu4����|��{Xmq��=�12������il��U2�u�3������`}�S��h�̜�O~�ww�U�<<==�B��o�M'Z�GW�Ԯ�i,d0����<�U�bI�;��/��^�W̶>%/�+?W����ɪ�ւ��r�3�)^�ڷ"����l��vh�3>��u���V'�n��D>�f��(�=-ii������<N��GʿD��O������?�2��Y^$�~n��Y��B�(�3SB�{�LG��J�jk}���P�	�sQ�������.4x��a����p��q�Q2��.zb�$�0�偣�
��~�K\�FP��JfLP�p��/ ��]J���{X3s�S�:5y����R�:e%�@9�I��뢏k?Z��r��ּ�#��^���Vר��ǻ��^w���|�;͘9�*=�f�P;�G)��7���j��$:�RL6Zx���1���~���]��/[��lBDo㬼k5��{ ��n���4Gd�A��Z��fB�~ZP�'�F�>�f��Z���:1���mZ5��R]��W�{#���R��/e��'<�z�j_o�����(
������Q���teUy#] '��xFZ���A׈o���X,%ʃ� �BDi��{3W��9�N�6/�ʘ�Ÿb�Ҝ�ꮦ���ν錑:# ��*������,}�sL,�:��jI�Ǌ�-)K(����j�{�w��H�G�I��R��O��_E���W��>�a
-���ڝ��Ţ��D!��dz׎|@0߇��ǻ:L�m�֜����x�(����K��V.�ͼ٬�a�5P��U(��텵nX�D���ʲ��w�r�Cф���w�|�?sm�ox6\j�[gV-��,��rϧ��3������g9�gG�������n��❯��
2��<&��[_@��jA�&�]z���+��οe=�~��*[�IE�6���G���Oť��CR�)�M>`�c���z���)o(��U�kX�Α,�	����ZPzR�O�W��]�e$�a]��2��i?!�`�B���Kw�.����i�"򢒖�ȥ\��M�D�b,k����[�������pv6Q^w��F:�Pm�����͛��Ͳ/כ��j�vuP͒g�]=A=���M���2��{|-���e-�$�"F0_����v��n��G�fd�`��ȝs�)�W��?�M��ǈ������PE۬��n`z����PY��s*4:W+�?��H�fh���A�|G��|��gع[�3З`(/�cv�f)c$X^�_Cm�G�3�$��Cfl�3�?�:�3'98�.�-wuO�.�R���˧�[�p�)[��C-�ѻү@P��ݨ46U��^�N��܄�H�DR��7�?y[,�kwI-��	�+���}�L�Vظ)�,KR �ԯ�Z8�{�k��+U��7�\��G�\Y8��'��������ri�n�x��0GJOc��cӱq9�K2�B(gW��s�WL���G�9`�g��كD�<��Yk�/j�����.�0{�QX�-�R�]�^����Q�L-��\	GO{H�u�="�`����싗�?����ED<�
0���;	&	.<�Dw�ʘ�)r��{�ccbՖm[9TtIA��kb�2n��J��IV�
x��Q
IG�ǩN���[���D~�����|�,�%X)K
��S��g���t��ȱ�o�4
@�i��x�z�ċ"
�ŰC���|F�o!�:�9`�=j/~���#J��M����BM��C���(s�����ڷw��� x�<��٬T�P�����󠓣#M�(�J�(@�����F+2���,!3�*�'[~:��g��������\��ğF�3��0=�-+�|�����*~���;�x;�jۜ�u��ޭJ��#Ck��&�Iީ�Jay�J�c� 3��h�
��P�c�:�g�nB�\����h�.���<��cUZXo�k�����,^�뵪�T|�4���A�7�̴�$c��rYj�fȓ��|Tz�g�	��t˛8r�6�!)gh���>{�{��\��L<�_�gth��Xc�Q��L������c�d����zf�$M�1t��g>��������"��6�����ZX�j�\S_�C����[]_�t8)c�>�0��)-���P��Ź|�&�*Z)B��Q����ҁ�As�ܱTl�g�ҡ��t;��NNOυv�b��"Y��q�(��RU��j-�<���ns�>����V�l�WEIQb���B�U}>i�F �T1pۨ�Z��Վz���)P�θ#���Q��9�����D�YJ+�M�inR�q&��u�fE��1�kv��A�n5���S LC�����8��L	���U��D��̔2�e�L��U}f	%BS�kD��'���P�{�_Dc�9ʹ��>�۟�g �[��GE��X��'o�Hڃ�����Z�%t�@�'nN	�vvq�L{"�U��듬)���A�EZ�(��c��~�N��I��a{��я~�Om�I�����-��2���n�.\�X����ל��ĭe����=�k���kr�S�1�RG�K��$��c��0����!�t!"��Lͫi�-����s��6�_�W�s1zlNOI���+��y5s�5'���՞ZE+����4��|�ݵ�{�<K�����N,q�6D'M�	¹��b�}��Uo���I���^���XmW���)]�N|1v�`�,d��`�V,[�Ӿό=:�v��1��Jb!,�)�74n�q�	������TI�!c��{�������4A\<�ύ���ԛ���ۺ����l�-����ۻ�k��}��i�@�RT�	,}���❦:Cܳ����	�`�\��G����!9KVG5:2����K��cϷ>��Oú�i)3�<���?��{�P^��e9�޴g�ؠd!O��á��mt+�ð�R�S䋚.#vX��_�ct�G���;v���|�u3�e�'���n�g��L�L�e N'�}䖂�o­�P�@t��"X��lH� �5�����L�����T  k&�M,綇H:��B\0�KK����6��7�K�t���!�ΜW4&�>�.IB��0�?B��'R���r��hoo4��W�D %_1��I1a\�e/D3�D+q4m�B����k��I�i�Ө�	`�}4P=��б� �]Sc��c�&��7i	Mf>�-P�9
����c����A{=�`�����fa�0��3��9�6n{GV����~z7��vb��)�+�H|��P|x^Ώ������r���M	�U�h���s/7�^��̧sK݉ie��,��9&c�A��fC�wxB��W�P����Yz���5�_"�՛�H�<U'�g��d����ʹA�Wމ����ᥢ�:M������u��v���>Agy)�z�����+��X�ĥR�M�[U�������a���Ӯ5kM��5��~7� An�rvp��� 5�U��HF�҃��CP٫Fn)�?_�"&����Y��>�k�"��]ˇ�g��I��䢹�7c��29��u��7�)�����l����:r������,��/~~�6P��ӳtl�`ƿ�5��R7���0������Ʈ�s0�p�����h���ſMMw/D�gh�a�V1�����vC9����fN��.�?(���C�q��YA ����8� ,X��A#.����{���m��9���}����
f�b��ݤR^Q8;f�8Z8VjA_AKc�7�C�e�W�Z�X}N��D�W�֊�9�g-ҧ�W�˹DKѓVb!��w�<�Ú�^���|F�$F��Y��V4�u�6�AF'v+�:�"����/�]>#�Tk�T��\����h%2�G�z��S���]��M���AI
��)گ�ǧ�1�L��Lw��S]��,[����=���1���zC&�Jp���a:��CsOv0˓�	ߝ��8�m��*����2��4'����Vn0N˫ �m�9��*ճ����k�HC���I�'.��ly!��C=��Ky���'La��j�M/.͘��`CYL9#Է8�T��wq)V_4�]�ŀر�3����=xA�{���pq#�������~o-�����B:]��(^�������������.K����@`N�s�k�����D.Ǉ�����[���8&��P��d��3L�'ٳS2�|G�\DW?�ړ��`as�����	4R�r:f���f���^���@�Cג3�Y�fC��H���e���R&��Ә(�c�WD��[�"�Fj��=h�/�f�d�Ku���J(�����<�(~`���걌�7��uǤs�Ԯ����0�1!�o����fx,��&y��ĺU�ȇwkd����2 �.،��3-�(�jXȻ�[�JI�n|��J�s`��;[Ӟ�P�u=�O{7����<a���FO��T#����:���󔫳����:#F�}jc ��/�GGO�*H����!��2ŋΡ >^IIovr���F	�ل���җ,��Є)h'��ݽˡ�����Y��-��������J������A�°�M��s�� Rp���6k�Pܑ�����F~��q��2���Wb�G��M�u�r �2BRI�mE�Ku�Pa�Ί��J@��������(C�ʊ\e�s#�b=��F�uc7�PF�����H��Nx��V)rKK/��rĻ�#�� ^�Ӈ��|��Cͯ�S��`g�2��U�8/�]ռ�b��^!�ח}k�0)�L�K��P���+���4Ýs�Љ�vz���Y���8��D7n�#YFhv��u5îR"i�fm%\!�6�[*�T�W�\�.��`s'�g����|�{������q�g����*Oʱ?e�b�W/IJ��X%����#P���F>~�)e��� l_����R�`$o�pZ;u	��?1�T˞R^�� p�>�͡4`�Gg�v�N�����ü@4g��2������]Oy1��z�J�]����cO��h���l�T��\S��H�Jd�e��� ]m�.����h4t���y4�Nt��B$�6���{!�����5z�3����A���Wq\�\�/�Wq����p�$�֨����t�~�L]CI���.�<9�d	����A���\�����nz���ۛ�[�w���:�贈K���f�p��a�v�3���S��}{���KaL���L��߅���A)�3/���r�ٕ�2;)i�R���}J���o�&�� jtz�2u��܂BL�?ϔ&Eܫ��@4톆��bA�Iu�̣E���4�»�����z���{ls����3؈�� 0}
�^O��q
�}�߭�Q�<����B�_%3�|�R��n˘��Z��r�gF��	+���Yw�7�����+�w����PK   �[SU;��I�Y  \  /   images/7842ad2d-d233-404b-8e7b-b5b626e67ff9.jpg��TM�.<X�� h��$�g��48�C�w h�������������s�9k�{���g�����ջ���v��U�<���W������ x^C� JK�����ʲ  �{I)Yd| ����$/E���E� � ��Of.N�����pG���4 �9���n�������_��w�6�p1 �����N�H9�������H�/���q���'�����p翍��/�)o�/���/?���pW��H;:y9[[}v����4w4����rq��w�:�9:;9:r�0�[����/���?=���D���v�_��}�7;��W�"�����?a����	�����?}d� j0  ��?u<� ����
�?uo�  �w @[��<@��������w�����/�^���&�#$$�#  "�|EDLAB@@FGFAEECCC���jJj�� �=�:..511��3�; H�H2(Ho �H(H�= ��mDEAB�/݃���Q0�0����H((�(hh�/0P�PQ��
* ��!�$:�� b�O�x���N)����ҁ	�'���U�<f.�2Z�]�x��uF��o��������D�W���������	����NC��Tb�(���kG&@! ���s�s#���7B���6l��&��_����]�Jp��."۪n�Xq*y��޸D�d8i�w�p�BG����_�+�s5Ү��H��oK�|��7�	ud<n%d�
���P���}�F�rV�*l�[D���l�����ۣ5���3 8x�Q14x<��^�Ѿ�i��Dz�ݻMũr"���^9.f�#̯>LD�/�yHk�h�;�df-'�O�����J8�����^G�y��F���5Ac��+�$��%Qא%F#֐��#��
�fH\�RÎ`�l��!��s�C��[M�����Ba�)J@�iuYN��~9Τ�9֘GA�fd[����K�B��3����;�]Ё�B~D����չ��f����NǲݣCJ~�ؖ�����5�R2CIӷ#�Ikyj
7v�	������Oލ�/Naq�c/C�A�R�2�g~\���avh��^ɷ�#
jq�T!1���U��W:�bƔ��Eͬ�I��K�� �]��y�F
q�	�q�!�z,��#�u����q}��{k�6�����=�5YU<�x�G�G�&=�V��ʪ��2Q>�j�	�� A�lu>$�/����|L^�T��λ�7�T��i������x����K�tr㞂��+P���P�ϓYL4a��xI��{O6ʥ:h��/�i�}���b��V_�S9�������� 
��"��U�_
�M[U�1��7��l7��w����]`���^��miQde��2�;pq=�p��7pj'V�pcQ>d�����<������M�n��ݫ=�u��[��-���1�����U�I�P��(	�Ө�N�-�~�m֏e�����S>�����1)_���x��X���_�~|�x���Cx^_|?'M�1�>����>�y
9�0�x���g�7X�yuy*����g���`0JR1(��h�������!3�,q�]0����Xa�\�3���>����!��W���Ũ�d|�Ѭ�H��&���dj�a}K�p?6�i�"4*OS7�YV�I�VX�>{�J�����U`�w�.~Ly}��U���ߐQ�"��>u=��q{�i>c0k��@-`����P��޵}�Av�ZҤg����(���X�~��ԡ�qE�����W���q������;�K^���`ھz�
��)8��2r�rs�tlEKV�<����쉗��Bm�[.,Rl�-�pD�d�U���� -+�W�����;gR|�[��vkWCˌ�?!߶������&II���0��ʥ7�l��Z��� aC�*��D�-�]��V1�i�~u`{�v�XW���d�T�:�PRK�fзؐ{������8� �N��I��q���=�!39�ؚ/�����vz��|W����<�=ed�W�5q(��)5����]1�
��!��s��Z9hD�*\�I��7�dp�����k3�q$�UMJDs��bߎ�%��Tl�g�����%̅7e�ٱj�OBYD��/����Pq��,�d��FZtH�^�;7?ǐ|����@ ��;٣�����;��D6�TG���� &q��L����b�(jJB��}#�yRkʣ�$R��Oڕqs
��@�/ku9,ƾ�f�_ǧ1_�,�oD�"|>h�Y?�1)Jr� �������T�����p�9����,G�t���?�-^7b�-�}_�T�5��c:T'���n*� �bZ3�D��b��[������|���x���L[#gc�Y}:}���_C_/y�m����tpas��I��oM����2	1��MZoOK3�`�)�Dw;d�O�E5�J\ה���*0o�v���	��,}?]"���(���W�����q��YP�5��c�]�QBl|qH�+�<�im�'��f�����I�?�W�ةW@1�I�e��JT@�5_��H�c�mL�ԏf��/>B� �����f^lRx�y�I�i��0[I,	�֮Ƣ�y,+�{��cb�����Q������w��L]do�>Z�o�7�AhU�6C��3�)�N�q�lQ�x��:a��3�Z�g�+n��W����x�x�4>'b�,�Qɛo�@_����)�ey"�-��y���N��^eIٲM���j�^۱���r�i�K�\Spp�o��ZEUί��2���/X3����b������u�V�u��x��}�&�1��4�\7�Y>n�v��|o1�Z�vֺ�!�x�T8�����7��{���
̈���?)�	!�zy>3е2� �9DL�x�l�V#�hX�2��\�*�4>A�=e�s��XLh��B� ���[�g ���ou���aƀ���	����`p�=?�gk:|�u=$Ȣ����ff�"X!h$N�>H�� 1�'X�|�C{D�%.}M���ӯ^���ʍ�C�N'�c��ՠ���>��.&=9��D~7Y��.6Z?�H{r�>�%�?��NBŴ1@��G(ا׬�c�*�Lh��PU!,X��kt98$=����_0��b�:��-�d|�?��d�h�#���%�����t���Y?��4���"�4��vb��@���Ԭ����!��A�f�4��z�I�|���ݸ���9�8/G<
�nF��|��kM��%Z_20���q_�X��b�:�۽Y-����g'���g+��)�>��܄v�iƭ�z�&��.f����(���a�vZ�l���4\TXKtZY@�}h#�K�2`�db]���dn,m������u�ӳjK[�:�f67�H2CU��ʳl�z�迌�����~;�v����a�$�w��eQԑ
C��%U� ���u�ǯ���
k�~tQ�vX��Y/���@��?���ʢ+RTAv񣪆����'K4�g4��	xsQ��+�)���V�jV���(
ڰ\0����Ǵc���7��Rn�M���~���IP?���h�'>�Î�f#9�l�N%:��u�]��o�{	�oc�%T����	�\TπS�mZppRN^.�:4ӳi�i����~a���2��%	[(]�����و�="9o�V�M��=�S�� ��"�ց-G��лӻM��t ��|1�^��+:�ׄb��y���o�Q���97�_��%_^��u�1�*�����O��YM����L�p�~�sL��SC�R^���Z�-U�K�d}��l���o���i*Y[�����AH��;%�ɇ��!�8Uo��,[C9��3_L'|��VA�P1ں�};����K�Sd��I�Q]���%���O�I �ߒW+�)�xN���@�,�*����l{R{�|vb��g�3���56��OZ0K�vX���z0���<�E�ãWv�YӒ�n�ےWkx��c�Wܒ�~��5sJx1���'��6;�/�ȵv�8��i�$��:��?�|~	�#�%�)<Q�y�B�-@8[������
�h�Q޲*9���ވtR��6��E�{;m;��r����e����h仈��O��v�AyT!KH���90"���0�d��A�G\���(���0��w.|�����-n@.�	Ҙ\��^|eC�t��K�|\��}%}��<�6+�s)}��%��*[g1��v�t�rH+Y��q-�	��||(	:d3h�K�u˧JG1���x�˽���'DE��/���LRp�F-W5��R+&$xlfh��[�֨�+�YEc&k����8�YMX�>7�s�+jdd�j��Wg[N��"�F��{|T�j�-!L���r���㈿UYR��L�`v�9a>��C,A�&�Y�37�m��\��%�qt���[���x�b��;MY�~d��P⪂xMN���;�O!V�X��np���]M���@/�KY}-�_ �+)K�k��&9���ﰷ�ZA{?����'q���98�C��X���5a\���I�m���w��i�W$�Į�2��v��!=1{�k=��h�ĵi�w�}���bc��t6ٌ5�Q�ظ�&ǫ�7���;lFm� �f{?����?����>i�I?h�"v��mYd�Y��_��4���li��H$FH�w�n��]k[{&���A�C�:�@.����xF�E��&�N��ܿ�S~+�#��T�g~=*0�_|��'Րc�ǵ%�d�4��\u.��e����;��7�1�v<D� �9B�	I���l�YT"&\U��j�3����S%v����f���D8m1E��b2��L���+ߗ4��@ة����Y��vCκٻ彾o8�5U�����֥j�SK�%o�IG�"�7w�HJ�!lW��G��mZ��V{ć�2 ��Lg;Y����exm:��|H�21��Bz٫�j/g�5�S	���(^�Ij-xL7�)����.��d<�]t���2�`f�|�V������#�>�x�~z��g\D	$�����L��I�+ʳ��4Mo��Pѐ���~f����6w$��
��տyo�a�	��
NN����(�6�S�� F^�`�d�?L�1ֿ���DP��4�ⲱ����v�h�����ۍ_��u�(��5�3t�i���#�^.*ų����M\��j�n���T�7AJ����m��A&�π����RqCw�7�Tr�5��W]�s�MÃMc�n�u�,�|/,:������p�Ƴ���;mO�඗��:��˺ߵ�7PwMK$W��mf-͐��k[х�b�|��u�5��7%����"P�#k0����Ak��q�o޾���s�������GJ��Q����`��~ls>�ga�����q�y��]�1N�/�w�&X�Ea!����vh�!F��~�O�U>���Q�r.G7:Z��|��bľ�՘�~O������A��c��V�*}oo�伮̱���]P��éV�m�}Y�f�'3��ZM�|���W�I�4��7>���_mf�0�X(�<��0�:C1�x����z�/?�P��A�@1j�K�$q�y�;]��.C��������j�g@��qW\����r��(��Ց�N�FW�[���D�n	7º��!!���8�%�j��-�|5�:�௽��`L��򋋂!@�&�M���/�S�}��(WN���Y���t�2��W��� ީ�!3�0�0{�\T�l�����Gxm�8��P(�)�/>#��u���[��Qt��-�T��	�L�+:�?h�fXl��GCmyjK�%��_���87��S��}�4>�7�� ��w��ܶ���?����g�S�(71��S��*5�)]z�b�F�ޙ�l������V��t�(�v_^R�r�]Q������n�T��%�(��<U�������,T�k�<�K�L,rC6��T���uV4��7���k�<F�j(�0�,�`N�I�&�h[�*n��R�!�D�&c�į���ʔ��m�H-���B��F�
��k;p��s����q���d�s���(�K�|�6Zl���������t&�^ɤ~ͺ�w�2�Hʴ�=隚�����NE�h��`{���||@�1�K.XrM_� �{��*}N�5�I�l��3����7�MF�]m�@�]��䞊I�/Ԭ��T���sBz=�"n I��9�1��o��(�׭!�����X��g�3/�B�O�&�W��	w\�cNmX�2(-���8��6�8��*c���ʏvo}���oq�1�����R@��gH�����YoHｼ�a�|�ήA���&�J�i�:]�Џ[�ܦg����4^�\��A�1�<��J���7�Wɥjp'�{�<)@W�i88t໗�8su/מ��u��	�:9�]�Ԟ4B��y0خ=��<�I)��^���@�Ӭ������tT���:A����h͹��S{��g�?rlHb�=\���]3МGF�Uv���T[.�\��@='J�����+���&���Ю��U1����7�"n�7��������F�TK�����.��3��#>A��ئ�ޚ��L:<�ݫ���UZ���Q�H6OP���0��1/��5��9�3ڣ�uMI����f[�h��r�h��u��Y��o/��&������/[������@L�\�{������R�Z0��(�#�ݔ��McbD�:�~�/�}�@x9x9�m<�g�R��.���[0�'ak�i�-9���9]���@��BɴwB�+�{~�0���N�+Db̐�����Yo�v]���0ډ��	�����&a���DU�s@��&���6~�/�6s(�#���g��G֙O	�X����V��c�_��xK�:V��b�Z(�c}.�
�<c��rw<��DڏTdH:�\�鳿W�%"���-���L����^a��_���Ǆo�b��g#�ڝ�E�B�J5���Nu�H���>:�ߞ��O�S	������jy'u�&�)�D�c��9:Dbѻ��K�,�\蝴rZ�>韒��	����\cZ�7�.��T8�l&x��/F}t��X2���P��K&��c��i�-�h�@L�:`E�$���璉���,uo���V%�Zۖ�"�s��ٮa����ɒ�`m�����z��Uc�c|_ΙԇX�����e����H��lmv�)\�H$� �j��5S۷�U��b�$p�̬���M����Ob_�B�EXg�8�½M$�c�J�Iĝ��TS�x�������Re�y����x�Z>�CI��J�z�9�iu�[���t*�O9�]���m�
kCu�z��{o�?Bz+��$E�맆iD[�'�g�Z����HZ��؊��}�9��|��^����Di|
�HF�u�r�n-rL���N�[�9��6!�Wq+.���x�3�)��S�[#���������Ao�,�w)�Z�!�1���`�=ےcp���^R
U7p	�S����i���S:�h|�~׆��S���I_za�I�Y���b�5#�+��C�����	z0��t���A�P�ꞦWaR���^�ox�Hț�P52uKI��({��`G�6mG�a��Z*�N�7�. �͢p&n4��Ն�$�q��SKZO�>U,�j��q3N�@!I􃶔���bK�'��>e=m[�y�����,����C�(Rj��az���:")$�/B�q2�f�W9E{��P��Ձa��K����C������D���Ɂ�U���~ۜ�[�����յThS��o���M+!oYp�}�jM&B��)���B��Lh�`����C�7j[3D�j!ޝ$r�8E�&�`���z�m�!2*^ANz��6����T�:�P�n�x�Sh؆���5���T/{K�F!��@�����ۯ;��h]{%������������U�E�{t�&��5za'�]�����9q@Ne�o��Ggŝ���	G�n*!z�z[?���C!�:-鵉�-P^5���n��@;�B�d]��^�Q��K[���Y��ϊd��vW!��Ӂ�|�����ϡɼ�"�Џ���m�A����R)�}��;�n.LzF{Z���@�M�9�@�1"���*�㺉A��ځ"�}�1�sx�
�����W4�����F(�)��d�������0����V�q��/�'���딽�.��Դx��AyL�񙥨��K��Q�uo1YP��~�oJv����(�cB���#���D����zb�PG(���@�PV�3 �����rV�P.�7�p=h$0��Sq(�z�MƗ䣮�3@~Q��g뇃�f�ж��
�#������m���[=�gPq�1N���yp��㤦]s5��f��~�ːߢ*�i����֠t��wgW���iޔK�j-���ߺ��g%�tkR�OB�ߏ�f\qp�2
I����<IL�5��&�+#-`'�x�Щ�o��o�h]?|wNykw���7t��%{#��\x�p�nt5Z���&��[�q�2a��A�U��۴`iX(
��� 7%yA���N�G�ӹ������P����x���m����s���_��l ��C��\��!aC��a���缯c��b��jo�-����ו�j����ȳrH{xj"�ݪ�á5����B2A׎���Yb(c�i�����	/�(9����~[ٜ$z*

�gc����~!���I{`�ļ
��㡤$��;�Ȳ>�q�!UOO
Oad4������v��v�p͹��Ҵm���bh͢n�P�!0�=H������I��mD����F�av�Rt�ϟI��<�[�z�9bY$��h!q]�������0i�(���BK��[��CH��z��\h�c��A�M�@�����LXT*�59:�?��L���j~܏ddv��o�L�raD=%�ŭS3�ОӺ�6�iߖ۟�{G;'!�~*�C�1��k�+�q��%]ݑ�z��z�������(�J������T�H=}�W�§��Bыg Vc,�5��w�&o���a�B�Am�Z��I�3]	�����SVC`$8�G-!`�+�����ӬjA(�3\��',#��7`{1ˏ'Q�Lf�����"wA�&ߚb0<�����3rV�ĸ�D_�ˁ!�<�,���b�S7��J	�' ��o��r+6��}`B�τO����ˏ-dM�o�9���2�E��F5�G�i��.��g�l���pb낀��ypg�G?0���~eݧH/�-����������l]ɸ=���[�du\)8�:�!��Vq<:�:S�F>k�_Q�������Ũ,�~B�j�=���H�՞���,�q���b�`Y��*�L�3�d���{`�g@����>�lR_?�#W�"@`�Wu�5=+e��O�Z=V���ˢ�����Vk���hec�RŘ��/x0�_E�479���	�RՉ�bX��,ӆ�Zt?>E7��%kl|��c�վ�^�ﻬ�{��ea�T�n�������L�T};f4����nɋmKF�����k!oZ꠾"�J;�D+����2uA�Ψ/]���e�j�����-��L��3hֿ��.�BطY���_����d���<����2��#m�k�������Rq���V����X���Z+S���� ���6�w��N%z�+�	�����О���P�L��dԣ^��,��e%/Qˡ��f��6��l���1�b�w�͒��s��)%�5���M�R�����M���� Դ���kD�e�ϾT�L<��Г�ԣrb{7A*��i����
9�3�[�{(^s��7�p�	.���8�1��܀�QvcS3Z�y��5+f
�~��s>�+B�g2Uy�}�+?�+�=)5�����8��?F�uy�k۴����Fe���[ڧ�G�~ZƆ�R�k�?��2 t�C.c�c�m�&�i�*0%eƅ͢��I.��<��Lۣeā� -퀨��^+�ڢr�Xs�o?*����iS�:���~5^s�t��!'?��Z�h�ʎ��!�QM��a��R�@�Q
7�{!�H
H����g���r�����.cⶈ�'Nl+�|P3�F���zB�T�:R�?�ݨdy+���)�
���%N�R�x��bl�^ٚ��F�cq�<x~^GG��O���Frz���p�=�@����b�3�˕��ZFŎ���4F�s$��du�Uk�br*������������ß7��
v�� ���á����S�2]�pVU��]��	�뎱t�G�~��ۃ7�%�3��gx�D�o	e��\��#ږ���?&�|GZb7�Գ.��D4���-�L���]�e��%A���I&#N��O4L�E�2���4���|��85�P��!3n�`i��E�)1Ih ���n�v���Q�q��2�ͨ��+���)��B�/N������� �j�kU�S�>� �[��������k��w�B�[�6,�xoDmK7��߅fN�I%m���r��7��)�`%�Q�=@5kbd� [d�ͼ6]^����Uk�b�v���qJ�f@�0��mv�6�,�qr��L�47�A��)��<!��Z��Q�z�iq��k�b2HT՘wQ�����
XHZ��Q���`��y/ 5�0�y��:���DcyW�z�������:���*%ú=��Yr�sX2UL@�(��J4��ɭ%ο�ι������Pi��u�#	N��g`Z�����Y�c`�)��B�	T�q~�ɵ�/����Hј���$�P����b�_g��>����Б5��p�p)Q.J�վ\����hq�p��ƏC��
�2
	�,��� Db-���;#qA�K�T+�[+#~�+͞Ǒh��zviv5���tcH*�#|<��w�E�C��x��^A�`�|ʘv,��FVe3]�� C�f����M��F��|Y�n���[gr�-"��/E�laE*�0hj����{�Z�o_�9��j���D#A�1f��.���M%w�r�����5��2�� �vc�Ⱥ��&�;a[��p�m�HS���B
�4+��[���������׋����_�S�|�ָ��<82*���j$�T
fQҸ�u
���*sk�
�I�X(����/&�;H��[pQ�ɑK)�S5o֢{�~���P�ů��չ!�r;��������p~��wh��P��j������8�q*��r�d������e����z���tvq�G�+$&��������(2�$Ϟܚ�q~���s{�����k�����ϼ� Y��k>F`�Gb�����6}n{&ςFCb����a¦�/غ��a�~|96�=S�#��~�_�vۆ�Z�o?g�Xܗق�Eꦆ���:O���ѽ��=������B	t0ou�>ya�����'ŕ[6�	,`�&Hy�U�T�*�
��i-d�L[@����}8�.��!B�$p�`s��	+����V5<:�휲0$����I�qei����F�4�vd�=Ⱦ�ۘx�!����]�*e��
귎*x�2��L*�4t�@`����ܨ�=Yj��Xԋ7F�;�%I�Ԇ������YAVu�g��w�5A�� ��X��I� ��:��M������@EP�q�����i�J(C�	�?�:<���KE����$C����[q�i0���h�X0�ʠ����;�$������{?:�K= +PD��lL�3��+C�����ئ���A��a�K�J��΃�U����"�����r	�a����ö���X�"u�Fo!�Ѡ����jrΦ{Nf�KP��7�euA{jN.�e����>wi��%�F��? C[ؕ���d=�Xt�" �"�.�p��}�=�7l'� 0K=`
(HW�R�/v^FM��튴Z æ+P� *�x����ݔ�����Ϧ8uYj�t�g8�Yg��
]DԤ�H<�^o�@M��,�FQ~ɓ�Mn�e���C��R@]�p^>)�<%��4J��f�@Q"l7Ue�<��`ؾ�*s0�3��ہE�o%N'������λ��^�:r��@>N:	P�<���I�G�g�� P���1�6�[ե�����?:��ߥAg�B�r#�����)0Rlã�e��Y����`B|W�N��)�<M��;T��ѝ�84`����(cz�L#�Mj���GTPc�]*̸9���̔�a�.��3�p��^ܲ�>A�ov���P�z'� ������4�fQcxCR��<�H�q�i�ď�m��:r�ɪ4��e�D�+�ͻ�q��@4���Ս��q5tZP[��.S�rM���#����b�u1���m�ná*�)��a,�J���챵
��"�=��r-�M�"��J�N���^Aɖ�g���I"A�/��,LcTx�4��NU]-��s�R�'M�]}� M�g � |�D���6�O��f�
�����KE�а��N���p���װ��|&��D:�9���۵�f�ȼ��� g(>���ݴ,z��d�����ŉ2 ����X��#e>)�����8�^(蓡���[+Sx��g�v 4������f�Ј!}� +�h�樽zƗ�"���f��jA��Nn�57��֏�5��_;J+�z �ky�䂘TB�H;���:�{غ��*��e�#~P����[��و�l���2C���sϳ_�����}�����2IZ9����Dw����].�<��#m�Ȓ��AP�]��m�q)�}��DM�?]�֜���|T,���Zx����]󱋨�@���״B�[I�Z�~�s]�����Y�!͟��F���z�W1p�5a����Cq���g~COR�k�(�f�W��_��&���첊!X��{O6��(Ȱ!ل�}��Q�l-#�a8p��
��v,d2�_R��(���>�Be;��bBN8�.k��ªѩ7�Ph��^�ugXAF��E��|�@�^�'6��x����
���㸋R�5�ѯ�
��D֝z�7.w�����[�-��@���a���ǝ�v������?�ep%�̒���"Ǻ2K������i�"�%��-n������O��j��1e~�,�C\���1��Ң�,�@|.�ܧ#���ݠ'���v~���G��b��K��H���a��n/��[��c�fY��&X��5�tF���՟��~U/��4�Q�F1Z_�4�l�P�&�W��7T4�/�Q�a���55AU`#A���b1�CHüe��Ơ���?Я��0'o��q/0U~�b�Mb����1�����ɛ���lR�� � ׺�A���V?�_=��8�P`@R�(��/��hj�W�P��4��1��×�.`˵�X���}�M�|��?�G�W	�k�R�?���)ݥI��qy|1���g >��l�����U�؈))���l�K�-�n��4wg���b�5���'��&7|�l�!����(kqg΢��h��]_���*�m�Ѳ���c`��`b����t��B�8Pٍ&�4�����~Ԃ�Ϧ���5�R�9�����ճu��S�f�U~���R�ؔˣ�F�����:6�	�KqNj����3���mɍ}�N�
��SW����e*�	�,��'��*��Af
j�?�}�^oQ$זsrHK�9S�4�;�w��Gz���L�O{�(���h��)��1+V���wi�?w��k?a��
do��.���>��:9��u�����ֈE���0����K����i�u�(�O'Np�/�rI��G"�孨���0,��6�I�6��L@+2^�ʦ��ƻ�ϊ.M5ѷ��1�
Ռ�M鈥U�5����h�z��]��y�A�t�x�6�Mk�|��_�0�.��'�`��E�h]ߴ&�d���o�:5}�� h(���J��X��T�qݎ��r�nԸ/5Ӭ=X_5��lm�ܧ�ZU[Tt�u����V����l��*���6K�0���,���ohedkj�]��_J<�Hz�Q0��_dLp�|{��:� Ny�QxM�:Ӌ�l��(��q_jⷰ��ER>�86�t�M�|��*��`3J>�?
[�.--�㭬�{/0-T����f\���:�U���"6d{IT��:��@�Y����Q�ǋ��z�ܤ�A�3����>v�r�G��X�/��o؜��^����_}�!���'@rV�1�r�;�=?A�N��#7g^"<��6��i����?���%b�#�2���ɂ�.��Ba�~�>��^�(Q /���m��	�L��dY@ʰ�ۅR��0�0^�&u�͍s��𓜴cb� (�A[e>j��w�����ߵ��Մ�t��RV���?�q%f��$�.�i��ph��#��4�f���۽-}���k�m��^��XF��Hbgʽ-�&����"6��2�/I��N�MV?ܔJ�W��!r��`����7f�qR�8�[ ���f���
��>��tL����W��4�fL����&�6�Z��Q��:Uw�l��f�7"�WhU��][#oc}�k�NYI�]��*�3��!��2�Yf�|'������S��q�P���|~���Cu�>Wr�OX�TV���n��� +�ݞ�s�+B7�����VBeQ۰�U#��<�y��T`��K>\`����w�AZF#�Ul��!���$`l���]`��=��r�9���z��RA��۟�m���1���(�lX��T�V�f}Q���^:,JX�;�l�i�"*��j��!���0B�!�=���cG$CG:��������"RN.3e;������#��k�t.n��D�4&�z�7���U'ӭ��(�*g�5͏l{���~䃴���]
ƭ�Q��m�殬���Ͽ��1�Р����G�WNSޖ� �/n߽h�5���'e,L���D��<�W�/�:�a��Ħ�6���
��/��5�"s�{�m:ײ�GyP���C��DMSƜ�K5"M�~5L�g ��x�Sї�񛹧���` �\��عlv�o��rBג$ەo�r�[����r�)[����)hONf�:6�Tx��c�k���8��xԵė�bMt�RR4��((��pL1v'�S�?i�����-��jo��Nl�����c��0Qi�85����=��+�CV'�þT��Z2	��^���o�]�Z�1�-%��r�	�N��Zʏs�a�g@��Q�������#nM��t
P�Z�����}��K
Z}2�H÷���rj�RQ�э�_��S� N�}���Y:���pJO���?2}֭�������y����tȑ��Uy5�N5)�D�M�\�t�M�3 ���
�qd��>�,tFF���_�����{�c�~�)  h�<=���������1L��$��bPCJ}��wگ����n�BNН �����ǺM����ŠU�khS9ql�3@R��3����̤�#�G�`����[�Lj�?�r�*(�Ѹ�}�p^��a��o$X <�!v�UO2|����t�Y2���1�a�FL�S:3�,[�ۤ5܎Z�%�$�%Zo(쎗���9����MC	���߮]*�dfI����{Ŕ��q�+����&Vg����Z�x��,c����2�WcE~��[�?DRUĪ9�z/!�n��k��|ҼƜ�e�\�d��~�C�N�a7#��k���Z˦���?B�s�X�oH#����0Ø&h�~�c5�m9*ј�r�^���s��q�_�eY��;��pa?J�-���M��R��@��6�[��J�\x�>�f��ϙ#K!��ʢ�/U/�Z�Λs�'z}\V����l�e���Z��Z� ����������$��By����A��L˳Iׯ��G����of�"����(��'�f��}+Mx�5����у��{���D��N��U����Ҝ��ջ>����4bvpU���	R2������v�z*��1��%�r�������yǖf]��%;��j[�`
���HQ��~����2����F��u��3��+�r�>%�1�Տ�`�(M>���1߇�S����]����-�7���l�y�,��o4���h>Jጨ�>ם/���q�čB�k��T��;���+�]�*�_�D2;O~����b*͉�����D��aك���� e]m9M��])��^?���8�l�+M�)�epI�ѻ��A�^�+H��E��c�U^��ŕG��r����҃v��C��Ӯ��*�!w͆� �[��oQ�5��5{��&�-��?�zw��7�ͻp!\!|¾���D��;%�4
J�q����
��DZ����)5��d�W2Y4!�:[n����t�׌ꤘw�m�ŋK!G��S��fEn��p�q�&s�
�s�����L�6�"`�^qT���CU�z����n1�*we-�����{�4���;\���{�'�*��	l��H%�w�G�K����������j���u(J� `��EZ �I��t!�����"�"$�H�  ���{�ޤIH�"���ͽg�s�w����k�^�5��p�2t�Af�(9��'F\�j�UЋ�������%�վA��G��4�{�dA�4�8�MXo9���|�z�r8�&X�D���V��q&��OG���[�1p׫.j�+�X���۷���%��BϚ�D>{'������q���Ñ%C��ؚ������SLUQD��}u�"[:1Ҽ���x�&m��H�ݓ
�O��])q��[r=P)<�@�=}�`�)d��K�h|<6�N���n�R卥�F7��
v<��k�	n�C�d�_w#�ݿ�"�)z�~&��.�����a����:�'���{˹�l=l�tu�j��H����w����:�|PC'w. o�_�L�~�!gS�	m��$z�H��FH�����%�(�@GҪ��_��}ri��ϟ� �6'�-z�磷dd�6�`bn}Э��|�?�]K���g��ɝ<o06����i��ɓl�'y�m�P����0 ���FA��t���d577h�V� <���E*��@����l{�V=�y|�{D���הL�M�oŏHD�oo���0���� �į�2+�V��4���9�B�D?�T�r�.�����Qï�F���D'E����ZS�-�iru%N����i�fv� OK�����ߴ�.�d<v�_mp��V	��Ƒ,�r+be��'�y=_�����[3���C���Ů=I�3ϭ/�2��$�K�	��Խ(k�UWf1��:M�����H4|7v�׃��C�ٴ]ד;Ǽ2d����*���	�:�b�&�����W�T�OL��d��{��+W�\���\�;l#Im��1�@�����<���B����F�.�^�f��j�&�$N�T�T{'���R�3�����3�.���F�p�I
�t���k���R�>p��	�9,��G89c~��(rCzb��Z�n�K�)��F�$� 11*ku[�FhJ��S�mY��to��p����^��/����z$Ί�?p^;�+���(��/X\��Mjo&I���V��W�%lAbI����W�j>����{B}to�g���zT@yh#C�e&L�Y�Q �GHp����܇'
e�Gs`��Ϭ ��bw�1������:�ڨ�IX��7)ۇ'� ��<uɃ��]�4�(=��;U:��ww>E<T�PA}� �	�t��U�Ȅ��?�U/ �Oׅ�RQ!�Vg~f.L��W�gO�Z��Ge�Ow�,�1�����6e0ό���p���$+_������|��;m����nc��&���p�����Γ�gx���>�g�S�꡸���Z�������mS����7��|9k��ڈ���w��,r�����ah�/4�ҡe��E�	�$�EDZ��La���1�dm�~��	�gd\�.^��Z)ǧ2�������[���~���o�'q�+�����.���
V�@�H�� ��@�N��);�0x�L"��oN��;���_j>AK��ͻ�Y����6-��:��.�=N1h2<.| ���?�7�����^�'k�I��!��WfO��,r�QJ,_�1Km�!���'�xb^��M�Z�Y��X�D��}b�1{;��n!j�O^^�Y�:+ �3e-���P���1խ��J�r8�$n��AC~�t�!�).�7"���\`�Q�0��<Y;g��������Ys�U�u�q��.�X;��a�q�2{�'���c�T�̅�<j����[L��v�)J���~��S��@ں �x��L��ضar��T'k����}-6��,��� �S�\�d7r��r�HJl�c�{Ӧ#�7Ĉ�x��./���э��LP��\��^bI)���\e�uN}A�.��r4+)4����Gv&��v�R=%vVk�*޳��$`�o�3��2�d8ۥG��\�͎q���!l:Yy*����?���F�y��{_<�Hv)��Eh���8�����h,A����K��J�	m�U|�FO��	l��&��k�A�A���Ś��L�7��QҞC���&K@�˕~���Xt\j6�eǓ��t:��NV d���<��ly�EG���9���׹�$4%�QA?7��P��ٯ�\g��&�z���3��ҿ�܄��x@�1�f6%0�76�����䭀T�g˂��矝�J=W� ���2�}*�Զ-k�݃Q�s	���59ш'l�� @E;B������/F���X�'���;D���>?-҆�:]�l%��3Gb��!��l< V^/�oe��Ȯ�O��>��Հ6#��\����'bj,�r/�q��9�}�^f�2޻��gf�n/�O)F4�X�%��-\�{�}��`������-��KN���K�U�1a8A��f�ӪK�x���4�T�&�K�� &�E�O/1���Gn��9}B����Ɨ0´�o�����{%�s���(+��^���O�=�RY�ӯj���a���FZ��l"sƴ-ޠ�2�rm��s�L�P�uk��� 0��~O�H+�~�����t��.��,!t��B�.N-u�I\I���t��#��!�@I���'Is��8�I��bB�7f���> ��e�WF=��Od��!�b�_)�����Is�n6�-�H��,r��yq78���|�����#��v�>cg���̯� o��a|3��p�:z��:-���4C߃Tqd����v��w=�l�܋�����Q`�ƫG�C�?����	m���2u9�_��&���ۿ�ebn��:���j18"�i�Uw:x�������3�	��x�
�{��. 3��-e����mEq�M6�f8��e�	�Y�����^�߸�Â�8�X����&�P8�.G�{�BM�}�u�xRO�V�#�7	�Z�-H�?������䝑-�������)l�(�~Y����d&�\+G�)��ݺ+�?M��,�׵�u(��ݾ�`]�O��0JW�G	���g�a|���-9�!��1㒝[���"��J����ؼ�N3{F����P�L��kⵜ���W��:B货4Im�2!��"�H����+��<�@\�>Al�uͮ��N���,�)k�d�Ώ�B��~d-5F�-
*�C���* �찢ꦻ��_T�F��]E_s^m�z��<k	�ě�\c��
O�(<�L:���G^��φ�+�/ ��ëk�tW�_�q��+�R3^0��Ul�$��d�Z�$�@Ѣ5]�o�����aj�%�\�~��h��a���%����h\�6��=m3�.w�TO�1q�Yõc�N�n�z.��9����l���W�S�gqK�*-�F�c��P�S4ts�%'�£5���g�F��j�f�5bf5Mhr�O��]s���,��� �Ѳ�3��-��YEH���	p�J�R�iApe[��<�<[����e��ʍe���6	M���8�u+Z�ޘ��%oQQ�y�筪	�?L1���QB;uBYA�Id�dC3R���@�������H���G-3@�]���T����.�_+�t���{��ki�?E��)y����*�3��S[>�W��`�c��g�|��n�T�j�D�Q�5C�򛄢��@��A�=���CN��v��- -���{��pN�$��zi�υ����t�?]Iǻ"��EE��sC+�O�M�"��]]�r���h=~���K �"�7wv�[��ݸ��s���'vø�L�J?�g�����z�"��Nߗ��u����?��
�%1'`n+�4�.�=L��s�SȞ&U�يT�Q�B��q�p���������e�T�xSߛУ+?<���(>�=�֐����8�G��w�`<��	SȽFY��g�讌��hL֗� h��6ˆf��#��*;�b��VFP	#HmDMw�Yu����H��b��A�A�F�G�*��+O��
-X�����������ʺ���`���,R���_�(���lv+G�R��/Hp�uK�۸&N��1��{^��l��F�dgP��~뻾�_�3���>5���}ҽ=@��U��r|�)QHA3�Z����+��T�L��n�*�$/\��d���8~��+�H��Yѐ��gopR�M��y��o[�8�&���8�cp7�^%�[q�lK�T�[,����yz9&&�Z�S��
��D�'�^���.W��i�A�o��8MY�m|Vn^o���e��d����+�~�C�Nj¢
��r��-sy��w��;T'�ү��Ȑ�	ء�#F�wV3{{��(??�7�`4]�N.n�pp䴗�7 �q�]	��A��uܸ��0ƿ���ѣ� �2b�5�G�Yj�i�j��ͩ���"Jwi��=	?X�U|�K��[�Gq��E�M�j�yj�[#k3B�GtC2�Ě�r���g�c�O�ء���AP��R�U�A���2�Kgc�������3;`��P��w��^7�S/����aI�Z�K�������L��@�"�==����*��G�@�>$�l���>��uļ��^1�7ϷU�������-�|��2��CAq3��#q&����ӡP>�Hs�vB!�l�@��x�!Ֆm/t���2-xX��f���۫E���<�l�/C{[C�tM���m��fK�/����',u���^�Bѩ�H�.
�I�cy����Q���CI�Z�&2i�Dq��l�&��ݾ��I�`]ܥz��`��aN|n�kr6��~���yG��/N%���M��HE�m}��!�j&^�jnZލ�ݷx��)Z$*�:�.d��ap���u.��z�^�Ɇ�ˑ�F�ܹ�,Vv;+�fG��]�&��{ӊ��܌
_�'�ats��9�J��_²��^����3���ԣ��������WK�M�����Q����Ň01�}���<���T�.w�튀�
2����)0�e��-��@=�.��H���?�.�j�hw^��:,��:z�ږƊ|n��*'�[s�r���c���9ٵZ��f`��jU�r 2���ĻVw�]��Z>-x��x=���V���(�%�_LfF���l�g0�z�̡C��8'5V3�Lu�f��GvRm�͔2z4�[^D��4
�-.b�Y�\�P���la�1�JY��50壈�&��S��v�!�4�O�cg��>���M���z�#��d���s�
�%���5��(!��5 R3-S��%��I�3��
hH���u�`����+�$��N��>���HW�s��d���F1���5���ƵǝCS�#g��~�೉I���*k[
�˵$� �tzj�h*��PE�m���'e�R�)_c��Oe����܍ "����2���(����z���O�ɥ�_'��A��+������~��=Z��������O��䧪/��f���
��ԩi����u@�'H��EI��`+�q����8+`Sa,!,H��u��Z�ZU�U�>-���wr=�\n��gM�*r�~v�_���Y!������9�9E���Є�_?17xV��`�N���YD�<���]=���:*Œf��=�V͹���QyD�F	_����H���P���j+p�sM����*����,`BAh��]��r�����c��C{Uvo�I����سB 
�%�v�截�i2�[PU�/�Z��z'K5�?��T�i2��.E���1�/�����-@�2�maH����E�Dك��X�''HB�`n�x��Yw�VV*�)/{�<�AS�_	�N�q�:	t4�g���)O&U�+��7�[]���xB ��`���\�@+� ��^�	��ˮX9�τjW��8nA7�t>��ʆ[Z�?��uV,`lO��f	>Gy�vU-{3JWW�#S:�I���� �� �1����GIm�_QRф).�iv{��h�ϫ��|HN�m���A[��AJa"G!����SlV�����==�"��Pt4Um~�+����y� ;�>�K���_l���6�3w��h�r�{�@a��a���C�)����P����=$�~t�1�Y�Ҁ��N�dr�vx�p��@����I>���p����u�Q��p�g�Ȗ�����i�K�ط����7ݿ+^/fD�6 ��M�M�8/�P�>T�@ad��$���P����::K�S�CN��TBD�y@��]C�D,��\����'��E_z��# ���8�W������;	�pbh��������+�Fd�sq{�:��S���PK   �[SU;��I�Y  \  /   images/943ec6f2-96cb-4ded-92cf-fc08d4cf4108.jpg��TM�.<X�� h��$�g��48�C�w h�������������s�9k�{���g�����ջ���v��U�<���W������ x^C� JK�����ʲ  �{I)Yd| ����$/E���E� � ��Of.N�����pG���4 �9���n�������_��w�6�p1 �����N�H9�������H�/���q���'�����p翍��/�)o�/���/?���pW��H;:y9[[}v����4w4����rq��w�:�9:;9:r�0�[����/���?=���D���v�_��}�7;��W�"�����?a����	�����?}d� j0  ��?u<� ����
�?uo�  �w @[��<@��������w�����/�^���&�#$$�#  "�|EDLAB@@FGFAEECCC���jJj�� �=�:..511��3�; H�H2(Ho �H(H�= ��mDEAB�/݃���Q0�0����H((�(hh�/0P�PQ��
* ��!�$:�� b�O�x���N)����ҁ	�'���U�<f.�2Z�]�x��uF��o��������D�W���������	����NC��Tb�(���kG&@! ���s�s#���7B���6l��&��_����]�Jp��."۪n�Xq*y��޸D�d8i�w�p�BG����_�+�s5Ү��H��oK�|��7�	ud<n%d�
���P���}�F�rV�*l�[D���l�����ۣ5���3 8x�Q14x<��^�Ѿ�i��Dz�ݻMũr"���^9.f�#̯>LD�/�yHk�h�;�df-'�O�����J8�����^G�y��F���5Ac��+�$��%Qא%F#֐��#��
�fH\�RÎ`�l��!��s�C��[M�����Ba�)J@�iuYN��~9Τ�9֘GA�fd[����K�B��3����;�]Ё�B~D����չ��f����NǲݣCJ~�ؖ�����5�R2CIӷ#�Ikyj
7v�	������Oލ�/Naq�c/C�A�R�2�g~\���avh��^ɷ�#
jq�T!1���U��W:�bƔ��Eͬ�I��K�� �]��y�F
q�	�q�!�z,��#�u����q}��{k�6�����=�5YU<�x�G�G�&=�V��ʪ��2Q>�j�	�� A�lu>$�/����|L^�T��λ�7�T��i������x����K�tr㞂��+P���P�ϓYL4a��xI��{O6ʥ:h��/�i�}���b��V_�S9�������� 
��"��U�_
�M[U�1��7��l7��w����]`���^��miQde��2�;pq=�p��7pj'V�pcQ>d�����<������M�n��ݫ=�u��[��-���1�����U�I�P��(	�Ө�N�-�~�m֏e�����S>�����1)_���x��X���_�~|�x���Cx^_|?'M�1�>����>�y
9�0�x���g�7X�yuy*����g���`0JR1(��h�������!3�,q�]0����Xa�\�3���>����!��W���Ũ�d|�Ѭ�H��&���dj�a}K�p?6�i�"4*OS7�YV�I�VX�>{�J�����U`�w�.~Ly}��U���ߐQ�"��>u=��q{�i>c0k��@-`����P��޵}�Av�ZҤg����(���X�~��ԡ�qE�����W���q������;�K^���`ھz�
��)8��2r�rs�tlEKV�<����쉗��Bm�[.,Rl�-�pD�d�U���� -+�W�����;gR|�[��vkWCˌ�?!߶������&II���0��ʥ7�l��Z��� aC�*��D�-�]��V1�i�~u`{�v�XW���d�T�:�PRK�fзؐ{������8� �N��I��q���=�!39�ؚ/�����vz��|W����<�=ed�W�5q(��)5����]1�
��!��s��Z9hD�*\�I��7�dp�����k3�q$�UMJDs��bߎ�%��Tl�g�����%̅7e�ٱj�OBYD��/����Pq��,�d��FZtH�^�;7?ǐ|����@ ��;٣�����;��D6�TG���� &q��L����b�(jJB��}#�yRkʣ�$R��Oڕqs
��@�/ku9,ƾ�f�_ǧ1_�,�oD�"|>h�Y?�1)Jr� �������T�����p�9����,G�t���?�-^7b�-�}_�T�5��c:T'���n*� �bZ3�D��b��[������|���x���L[#gc�Y}:}���_C_/y�m����tpas��I��oM����2	1��MZoOK3�`�)�Dw;d�O�E5�J\ה���*0o�v���	��,}?]"���(���W�����q��YP�5��c�]�QBl|qH�+�<�im�'��f�����I�?�W�ةW@1�I�e��JT@�5_��H�c�mL�ԏf��/>B� �����f^lRx�y�I�i��0[I,	�֮Ƣ�y,+�{��cb�����Q������w��L]do�>Z�o�7�AhU�6C��3�)�N�q�lQ�x��:a��3�Z�g�+n��W����x�x�4>'b�,�Qɛo�@_����)�ey"�-��y���N��^eIٲM���j�^۱���r�i�K�\Spp�o��ZEUί��2���/X3����b������u�V�u��x��}�&�1��4�\7�Y>n�v��|o1�Z�vֺ�!�x�T8�����7��{���
̈���?)�	!�zy>3е2� �9DL�x�l�V#�hX�2��\�*�4>A�=e�s��XLh��B� ���[�g ���ou���aƀ���	����`p�=?�gk:|�u=$Ȣ����ff�"X!h$N�>H�� 1�'X�|�C{D�%.}M���ӯ^���ʍ�C�N'�c��ՠ���>��.&=9��D~7Y��.6Z?�H{r�>�%�?��NBŴ1@��G(ا׬�c�*�Lh��PU!,X��kt98$=����_0��b�:��-�d|�?��d�h�#���%�����t���Y?��4���"�4��vb��@���Ԭ����!��A�f�4��z�I�|���ݸ���9�8/G<
�nF��|��kM��%Z_20���q_�X��b�:�۽Y-����g'���g+��)�>��܄v�iƭ�z�&��.f����(���a�vZ�l���4\TXKtZY@�}h#�K�2`�db]���dn,m������u�ӳjK[�:�f67�H2CU��ʳl�z�迌�����~;�v����a�$�w��eQԑ
C��%U� ���u�ǯ���
k�~tQ�vX��Y/���@��?���ʢ+RTAv񣪆����'K4�g4��	xsQ��+�)���V�jV���(
ڰ\0����Ǵc���7��Rn�M���~���IP?���h�'>�Î�f#9�l�N%:��u�]��o�{	�oc�%T����	�\TπS�mZppRN^.�:4ӳi�i����~a���2��%	[(]�����و�="9o�V�M��=�S�� ��"�ց-G��лӻM��t ��|1�^��+:�ׄb��y���o�Q���97�_��%_^��u�1�*�����O��YM����L�p�~�sL��SC�R^���Z�-U�K�d}��l���o���i*Y[�����AH��;%�ɇ��!�8Uo��,[C9��3_L'|��VA�P1ں�};����K�Sd��I�Q]���%���O�I �ߒW+�)�xN���@�,�*����l{R{�|vb��g�3���56��OZ0K�vX���z0���<�E�ãWv�YӒ�n�ےWkx��c�Wܒ�~��5sJx1���'��6;�/�ȵv�8��i�$��:��?�|~	�#�%�)<Q�y�B�-@8[������
�h�Q޲*9���ވtR��6��E�{;m;��r����e����h仈��O��v�AyT!KH���90"���0�d��A�G\���(���0��w.|�����-n@.�	Ҙ\��^|eC�t��K�|\��}%}��<�6+�s)}��%��*[g1��v�t�rH+Y��q-�	��||(	:d3h�K�u˧JG1���x�˽���'DE��/���LRp�F-W5��R+&$xlfh��[�֨�+�YEc&k����8�YMX�>7�s�+jdd�j��Wg[N��"�F��{|T�j�-!L���r���㈿UYR��L�`v�9a>��C,A�&�Y�37�m��\��%�qt���[���x�b��;MY�~d��P⪂xMN���;�O!V�X��np���]M���@/�KY}-�_ �+)K�k��&9���ﰷ�ZA{?����'q���98�C��X���5a\���I�m���w��i�W$�Į�2��v��!=1{�k=��h�ĵi�w�}���bc��t6ٌ5�Q�ظ�&ǫ�7���;lFm� �f{?����?����>i�I?h�"v��mYd�Y��_��4���li��H$FH�w�n��]k[{&���A�C�:�@.����xF�E��&�N��ܿ�S~+�#��T�g~=*0�_|��'Րc�ǵ%�d�4��\u.��e����;��7�1�v<D� �9B�	I���l�YT"&\U��j�3����S%v����f���D8m1E��b2��L���+ߗ4��@ة����Y��vCκٻ彾o8�5U�����֥j�SK�%o�IG�"�7w�HJ�!lW��G��mZ��V{ć�2 ��Lg;Y����exm:��|H�21��Bz٫�j/g�5�S	���(^�Ij-xL7�)����.��d<�]t���2�`f�|�V������#�>�x�~z��g\D	$�����L��I�+ʳ��4Mo��Pѐ���~f����6w$��
��տyo�a�	��
NN����(�6�S�� F^�`�d�?L�1ֿ���DP��4�ⲱ����v�h�����ۍ_��u�(��5�3t�i���#�^.*ų����M\��j�n���T�7AJ����m��A&�π����RqCw�7�Tr�5��W]�s�MÃMc�n�u�,�|/,:������p�Ƴ���;mO�඗��:��˺ߵ�7PwMK$W��mf-͐��k[х�b�|��u�5��7%����"P�#k0����Ak��q�o޾���s�������GJ��Q����`��~ls>�ga�����q�y��]�1N�/�w�&X�Ea!����vh�!F��~�O�U>���Q�r.G7:Z��|��bľ�՘�~O������A��c��V�*}oo�伮̱���]P��éV�m�}Y�f�'3��ZM�|���W�I�4��7>���_mf�0�X(�<��0�:C1�x����z�/?�P��A�@1j�K�$q�y�;]��.C��������j�g@��qW\����r��(��Ց�N�FW�[���D�n	7º��!!���8�%�j��-�|5�:�௽��`L��򋋂!@�&�M���/�S�}��(WN���Y���t�2��W��� ީ�!3�0�0{�\T�l�����Gxm�8��P(�)�/>#��u���[��Qt��-�T��	�L�+:�?h�fXl��GCmyjK�%��_���87��S��}�4>�7�� ��w��ܶ���?����g�S�(71��S��*5�)]z�b�F�ޙ�l������V��t�(�v_^R�r�]Q������n�T��%�(��<U�������,T�k�<�K�L,rC6��T���uV4��7���k�<F�j(�0�,�`N�I�&�h[�*n��R�!�D�&c�į���ʔ��m�H-���B��F�
��k;p��s����q���d�s���(�K�|�6Zl���������t&�^ɤ~ͺ�w�2�Hʴ�=隚�����NE�h��`{���||@�1�K.XrM_� �{��*}N�5�I�l��3����7�MF�]m�@�]��䞊I�/Ԭ��T���sBz=�"n I��9�1��o��(�׭!�����X��g�3/�B�O�&�W��	w\�cNmX�2(-���8��6�8��*c���ʏvo}���oq�1�����R@��gH�����YoHｼ�a�|�ήA���&�J�i�:]�Џ[�ܦg����4^�\��A�1�<��J���7�Wɥjp'�{�<)@W�i88t໗�8su/מ��u��	�:9�]�Ԟ4B��y0خ=��<�I)��^���@�Ӭ������tT���:A����h͹��S{��g�?rlHb�=\���]3МGF�Uv���T[.�\��@='J�����+���&���Ю��U1����7�"n�7��������F�TK�����.��3��#>A��ئ�ޚ��L:<�ݫ���UZ���Q�H6OP���0��1/��5��9�3ڣ�uMI����f[�h��r�h��u��Y��o/��&������/[������@L�\�{������R�Z0��(�#�ݔ��McbD�:�~�/�}�@x9x9�m<�g�R��.���[0�'ak�i�-9���9]���@��BɴwB�+�{~�0���N�+Db̐�����Yo�v]���0ډ��	�����&a���DU�s@��&���6~�/�6s(�#���g��G֙O	�X����V��c�_��xK�:V��b�Z(�c}.�
�<c��rw<��DڏTdH:�\�鳿W�%"���-���L����^a��_���Ǆo�b��g#�ڝ�E�B�J5���Nu�H���>:�ߞ��O�S	������jy'u�&�)�D�c��9:Dbѻ��K�,�\蝴rZ�>韒��	����\cZ�7�.��T8�l&x��/F}t��X2���P��K&��c��i�-�h�@L�:`E�$���璉���,uo���V%�Zۖ�"�s��ٮa����ɒ�`m�����z��Uc�c|_ΙԇX�����e����H��lmv�)\�H$� �j��5S۷�U��b�$p�̬���M����Ob_�B�EXg�8�½M$�c�J�Iĝ��TS�x�������Re�y����x�Z>�CI��J�z�9�iu�[���t*�O9�]���m�
kCu�z��{o�?Bz+��$E�맆iD[�'�g�Z����HZ��؊��}�9��|��^����Di|
�HF�u�r�n-rL���N�[�9��6!�Wq+.���x�3�)��S�[#���������Ao�,�w)�Z�!�1���`�=ےcp���^R
U7p	�S����i���S:�h|�~׆��S���I_za�I�Y���b�5#�+��C�����	z0��t���A�P�ꞦWaR���^�ox�Hț�P52uKI��({��`G�6mG�a��Z*�N�7�. �͢p&n4��Ն�$�q��SKZO�>U,�j��q3N�@!I􃶔���bK�'��>e=m[�y�����,����C�(Rj��az���:")$�/B�q2�f�W9E{��P��Ձa��K����C������D���Ɂ�U���~ۜ�[�����յThS��o���M+!oYp�}�jM&B��)���B��Lh�`����C�7j[3D�j!ޝ$r�8E�&�`���z�m�!2*^ANz��6����T�:�P�n�x�Sh؆���5���T/{K�F!��@�����ۯ;��h]{%������������U�E�{t�&��5za'�]�����9q@Ne�o��Ggŝ���	G�n*!z�z[?���C!�:-鵉�-P^5���n��@;�B�d]��^�Q��K[���Y��ϊd��vW!��Ӂ�|�����ϡɼ�"�Џ���m�A����R)�}��;�n.LzF{Z���@�M�9�@�1"���*�㺉A��ځ"�}�1�sx�
�����W4�����F(�)��d�������0����V�q��/�'���딽�.��Դx��AyL�񙥨��K��Q�uo1YP��~�oJv����(�cB���#���D����zb�PG(���@�PV�3 �����rV�P.�7�p=h$0��Sq(�z�MƗ䣮�3@~Q��g뇃�f�ж��
�#������m���[=�gPq�1N���yp��㤦]s5��f��~�ːߢ*�i����֠t��wgW���iޔK�j-���ߺ��g%�tkR�OB�ߏ�f\qp�2
I����<IL�5��&�+#-`'�x�Щ�o��o�h]?|wNykw���7t��%{#��\x�p�nt5Z���&��[�q�2a��A�U��۴`iX(
��� 7%yA���N�G�ӹ������P����x���m����s���_��l ��C��\��!aC��a���缯c��b��jo�-����ו�j����ȳrH{xj"�ݪ�á5����B2A׎���Yb(c�i�����	/�(9����~[ٜ$z*

�gc����~!���I{`�ļ
��㡤$��;�Ȳ>�q�!UOO
Oad4������v��v�p͹��Ҵm���bh͢n�P�!0�=H������I��mD����F�av�Rt�ϟI��<�[�z�9bY$��h!q]�������0i�(���BK��[��CH��z��\h�c��A�M�@�����LXT*�59:�?��L���j~܏ddv��o�L�raD=%�ŭS3�ОӺ�6�iߖ۟�{G;'!�~*�C�1��k�+�q��%]ݑ�z��z�������(�J������T�H=}�W�§��Bыg Vc,�5��w�&o���a�B�Am�Z��I�3]	�����SVC`$8�G-!`�+�����ӬjA(�3\��',#��7`{1ˏ'Q�Lf�����"wA�&ߚb0<�����3rV�ĸ�D_�ˁ!�<�,���b�S7��J	�' ��o��r+6��}`B�τO����ˏ-dM�o�9���2�E��F5�G�i��.��g�l���pb낀��ypg�G?0���~eݧH/�-����������l]ɸ=���[�du\)8�:�!��Vq<:�:S�F>k�_Q�������Ũ,�~B�j�=���H�՞���,�q���b�`Y��*�L�3�d���{`�g@����>�lR_?�#W�"@`�Wu�5=+e��O�Z=V���ˢ�����Vk���hec�RŘ��/x0�_E�479���	�RՉ�bX��,ӆ�Zt?>E7��%kl|��c�վ�^�ﻬ�{��ea�T�n�������L�T};f4����nɋmKF�����k!oZ꠾"�J;�D+����2uA�Ψ/]���e�j�����-��L��3hֿ��.�BطY���_����d���<����2��#m�k�������Rq���V����X���Z+S���� ���6�w��N%z�+�	�����О���P�L��dԣ^��,��e%/Qˡ��f��6��l���1�b�w�͒��s��)%�5���M�R�����M���� Դ���kD�e�ϾT�L<��Г�ԣrb{7A*��i����
9�3�[�{(^s��7�p�	.���8�1��܀�QvcS3Z�y��5+f
�~��s>�+B�g2Uy�}�+?�+�=)5�����8��?F�uy�k۴����Fe���[ڧ�G�~ZƆ�R�k�?��2 t�C.c�c�m�&�i�*0%eƅ͢��I.��<��Lۣeā� -퀨��^+�ڢr�Xs�o?*����iS�:���~5^s�t��!'?��Z�h�ʎ��!�QM��a��R�@�Q
7�{!�H
H����g���r�����.cⶈ�'Nl+�|P3�F���zB�T�:R�?�ݨdy+���)�
���%N�R�x��bl�^ٚ��F�cq�<x~^GG��O���Frz���p�=�@����b�3�˕��ZFŎ���4F�s$��du�Uk�br*������������ß7��
v�� ���á����S�2]�pVU��]��	�뎱t�G�~��ۃ7�%�3��gx�D�o	e��\��#ږ���?&�|GZb7�Գ.��D4���-�L���]�e��%A���I&#N��O4L�E�2���4���|��85�P��!3n�`i��E�)1Ih ���n�v���Q�q��2�ͨ��+���)��B�/N������� �j�kU�S�>� �[��������k��w�B�[�6,�xoDmK7��߅fN�I%m���r��7��)�`%�Q�=@5kbd� [d�ͼ6]^����Uk�b�v���qJ�f@�0��mv�6�,�qr��L�47�A��)��<!��Z��Q�z�iq��k�b2HT՘wQ�����
XHZ��Q���`��y/ 5�0�y��:���DcyW�z�������:���*%ú=��Yr�sX2UL@�(��J4��ɭ%ο�ι������Pi��u�#	N��g`Z�����Y�c`�)��B�	T�q~�ɵ�/����Hј���$�P����b�_g��>����Б5��p�p)Q.J�վ\����hq�p��ƏC��
�2
	�,��� Db-���;#qA�K�T+�[+#~�+͞Ǒh��zviv5���tcH*�#|<��w�E�C��x��^A�`�|ʘv,��FVe3]�� C�f����M��F��|Y�n���[gr�-"��/E�laE*�0hj����{�Z�o_�9��j���D#A�1f��.���M%w�r�����5��2�� �vc�Ⱥ��&�;a[��p�m�HS���B
�4+��[���������׋����_�S�|�ָ��<82*���j$�T
fQҸ�u
���*sk�
�I�X(����/&�;H��[pQ�ɑK)�S5o֢{�~���P�ů��չ!�r;��������p~��wh��P��j������8�q*��r�d������e����z���tvq�G�+$&��������(2�$Ϟܚ�q~���s{�����k�����ϼ� Y��k>F`�Gb�����6}n{&ςFCb����a¦�/غ��a�~|96�=S�#��~�_�vۆ�Z�o?g�Xܗق�Eꦆ���:O���ѽ��=������B	t0ou�>ya�����'ŕ[6�	,`�&Hy�U�T�*�
��i-d�L[@����}8�.��!B�$p�`s��	+����V5<:�휲0$����I�qei����F�4�vd�=Ⱦ�ۘx�!����]�*e��
귎*x�2��L*�4t�@`����ܨ�=Yj��Xԋ7F�;�%I�Ԇ������YAVu�g��w�5A�� ��X��I� ��:��M������@EP�q�����i�J(C�	�?�:<���KE����$C����[q�i0���h�X0�ʠ����;�$������{?:�K= +PD��lL�3��+C�����ئ���A��a�K�J��΃�U����"�����r	�a����ö���X�"u�Fo!�Ѡ����jrΦ{Nf�KP��7�euA{jN.�e����>wi��%�F��? C[ؕ���d=�Xt�" �"�.�p��}�=�7l'� 0K=`
(HW�R�/v^FM��튴Z æ+P� *�x����ݔ�����Ϧ8uYj�t�g8�Yg��
]DԤ�H<�^o�@M��,�FQ~ɓ�Mn�e���C��R@]�p^>)�<%��4J��f�@Q"l7Ue�<��`ؾ�*s0�3��ہE�o%N'������λ��^�:r��@>N:	P�<���I�G�g�� P���1�6�[ե�����?:��ߥAg�B�r#�����)0Rlã�e��Y����`B|W�N��)�<M��;T��ѝ�84`����(cz�L#�Mj���GTPc�]*̸9���̔�a�.��3�p��^ܲ�>A�ov���P�z'� ������4�fQcxCR��<�H�q�i�ď�m��:r�ɪ4��e�D�+�ͻ�q��@4���Ս��q5tZP[��.S�rM���#����b�u1���m�ná*�)��a,�J���챵
��"�=��r-�M�"��J�N���^Aɖ�g���I"A�/��,LcTx�4��NU]-��s�R�'M�]}� M�g � |�D���6�O��f�
�����KE�а��N���p���װ��|&��D:�9���۵�f�ȼ��� g(>���ݴ,z��d�����ŉ2 ����X��#e>)�����8�^(蓡���[+Sx��g�v 4������f�Ј!}� +�h�樽zƗ�"���f��jA��Nn�57��֏�5��_;J+�z �ky�䂘TB�H;���:�{غ��*��e�#~P����[��و�l���2C���sϳ_�����}�����2IZ9����Dw����].�<��#m�Ȓ��AP�]��m�q)�}��DM�?]�֜���|T,���Zx����]󱋨�@���״B�[I�Z�~�s]�����Y�!͟��F���z�W1p�5a����Cq���g~COR�k�(�f�W��_��&���첊!X��{O6��(Ȱ!ل�}��Q�l-#�a8p��
��v,d2�_R��(���>�Be;��bBN8�.k��ªѩ7�Ph��^�ugXAF��E��|�@�^�'6��x����
���㸋R�5�ѯ�
��D֝z�7.w�����[�-��@���a���ǝ�v������?�ep%�̒���"Ǻ2K������i�"�%��-n������O��j��1e~�,�C\���1��Ң�,�@|.�ܧ#���ݠ'���v~���G��b��K��H���a��n/��[��c�fY��&X��5�tF���՟��~U/��4�Q�F1Z_�4�l�P�&�W��7T4�/�Q�a���55AU`#A���b1�CHüe��Ơ���?Я��0'o��q/0U~�b�Mb����1�����ɛ���lR�� � ׺�A���V?�_=��8�P`@R�(��/��hj�W�P��4��1��×�.`˵�X���}�M�|��?�G�W	�k�R�?���)ݥI��qy|1���g >��l�����U�؈))���l�K�-�n��4wg���b�5���'��&7|�l�!����(kqg΢��h��]_���*�m�Ѳ���c`��`b����t��B�8Pٍ&�4�����~Ԃ�Ϧ���5�R�9�����ճu��S�f�U~���R�ؔˣ�F�����:6�	�KqNj����3���mɍ}�N�
��SW����e*�	�,��'��*��Af
j�?�}�^oQ$זsrHK�9S�4�;�w��Gz���L�O{�(���h��)��1+V���wi�?w��k?a��
do��.���>��:9��u�����ֈE���0����K����i�u�(�O'Np�/�rI��G"�孨���0,��6�I�6��L@+2^�ʦ��ƻ�ϊ.M5ѷ��1�
Ռ�M鈥U�5����h�z��]��y�A�t�x�6�Mk�|��_�0�.��'�`��E�h]ߴ&�d���o�:5}�� h(���J��X��T�qݎ��r�nԸ/5Ӭ=X_5��lm�ܧ�ZU[Tt�u����V����l��*���6K�0���,���ohedkj�]��_J<�Hz�Q0��_dLp�|{��:� Ny�QxM�:Ӌ�l��(��q_jⷰ��ER>�86�t�M�|��*��`3J>�?
[�.--�㭬�{/0-T����f\���:�U���"6d{IT��:��@�Y����Q�ǋ��z�ܤ�A�3����>v�r�G��X�/��o؜��^����_}�!���'@rV�1�r�;�=?A�N��#7g^"<��6��i����?���%b�#�2���ɂ�.��Ba�~�>��^�(Q /���m��	�L��dY@ʰ�ۅR��0�0^�&u�͍s��𓜴cb� (�A[e>j��w�����ߵ��Մ�t��RV���?�q%f��$�.�i��ph��#��4�f���۽-}���k�m��^��XF��Hbgʽ-�&����"6��2�/I��N�MV?ܔJ�W��!r��`����7f�qR�8�[ ���f���
��>��tL����W��4�fL����&�6�Z��Q��:Uw�l��f�7"�WhU��][#oc}�k�NYI�]��*�3��!��2�Yf�|'������S��q�P���|~���Cu�>Wr�OX�TV���n��� +�ݞ�s�+B7�����VBeQ۰�U#��<�y��T`��K>\`����w�AZF#�Ul��!���$`l���]`��=��r�9���z��RA��۟�m���1���(�lX��T�V�f}Q���^:,JX�;�l�i�"*��j��!���0B�!�=���cG$CG:��������"RN.3e;������#��k�t.n��D�4&�z�7���U'ӭ��(�*g�5͏l{���~䃴���]
ƭ�Q��m�殬���Ͽ��1�Р����G�WNSޖ� �/n߽h�5���'e,L���D��<�W�/�:�a��Ħ�6���
��/��5�"s�{�m:ײ�GyP���C��DMSƜ�K5"M�~5L�g ��x�Sї�񛹧���` �\��عlv�o��rBג$ەo�r�[����r�)[����)hONf�:6�Tx��c�k���8��xԵė�bMt�RR4��((��pL1v'�S�?i�����-��jo��Nl�����c��0Qi�85����=��+�CV'�þT��Z2	��^���o�]�Z�1�-%��r�	�N��Zʏs�a�g@��Q�������#nM��t
P�Z�����}��K
Z}2�H÷���rj�RQ�э�_��S� N�}���Y:���pJO���?2}֭�������y����tȑ��Uy5�N5)�D�M�\�t�M�3 ���
�qd��>�,tFF���_�����{�c�~�)  h�<=���������1L��$��bPCJ}��wگ����n�BNН �����ǺM����ŠU�khS9ql�3@R��3����̤�#�G�`����[�Lj�?�r�*(�Ѹ�}�p^��a��o$X <�!v�UO2|����t�Y2���1�a�FL�S:3�,[�ۤ5܎Z�%�$�%Zo(쎗���9����MC	���߮]*�dfI����{Ŕ��q�+����&Vg����Z�x��,c����2�WcE~��[�?DRUĪ9�z/!�n��k��|ҼƜ�e�\�d��~�C�N�a7#��k���Z˦���?B�s�X�oH#����0Ø&h�~�c5�m9*ј�r�^���s��q�_�eY��;��pa?J�-���M��R��@��6�[��J�\x�>�f��ϙ#K!��ʢ�/U/�Z�Λs�'z}\V����l�e���Z��Z� ����������$��By����A��L˳Iׯ��G����of�"����(��'�f��}+Mx�5����у��{���D��N��U����Ҝ��ջ>����4bvpU���	R2������v�z*��1��%�r�������yǖf]��%;��j[�`
���HQ��~����2����F��u��3��+�r�>%�1�Տ�`�(M>���1߇�S����]����-�7���l�y�,��o4���h>Jጨ�>ם/���q�čB�k��T��;���+�]�*�_�D2;O~����b*͉�����D��aك���� e]m9M��])��^?���8�l�+M�)�epI�ѻ��A�^�+H��E��c�U^��ŕG��r����҃v��C��Ӯ��*�!w͆� �[��oQ�5��5{��&�-��?�zw��7�ͻp!\!|¾���D��;%�4
J�q����
��DZ����)5��d�W2Y4!�:[n����t�׌ꤘw�m�ŋK!G��S��fEn��p�q�&s�
�s�����L�6�"`�^qT���CU�z����n1�*we-�����{�4���;\���{�'�*��	l��H%�w�G�K����������j���u(J� `��EZ �I��t!�����"�"$�H�  ���{�ޤIH�"���ͽg�s�w����k�^�5��p�2t�Af�(9��'F\�j�UЋ�������%�վA��G��4�{�dA�4�8�MXo9���|�z�r8�&X�D���V��q&��OG���[�1p׫.j�+�X���۷���%��BϚ�D>{'������q���Ñ%C��ؚ������SLUQD��}u�"[:1Ҽ���x�&m��H�ݓ
�O��])q��[r=P)<�@�=}�`�)d��K�h|<6�N���n�R卥�F7��
v<��k�	n�C�d�_w#�ݿ�"�)z�~&��.�����a����:�'���{˹�l=l�tu�j��H����w����:�|PC'w. o�_�L�~�!gS�	m��$z�H��FH�����%�(�@GҪ��_��}ri��ϟ� �6'�-z�磷dd�6�`bn}Э��|�?�]K���g��ɝ<o06����i��ɓl�'y�m�P����0 ���FA��t���d577h�V� <���E*��@����l{�V=�y|�{D���הL�M�oŏHD�oo���0���� �į�2+�V��4���9�B�D?�T�r�.�����Qï�F���D'E����ZS�-�iru%N����i�fv� OK�����ߴ�.�d<v�_mp��V	��Ƒ,�r+be��'�y=_�����[3���C���Ů=I�3ϭ/�2��$�K�	��Խ(k�UWf1��:M�����H4|7v�׃��C�ٴ]ד;Ǽ2d����*���	�:�b�&�����W�T�OL��d��{��+W�\���\�;l#Im��1�@�����<���B����F�.�^�f��j�&�$N�T�T{'���R�3�����3�.���F�p�I
�t���k���R�>p��	�9,��G89c~��(rCzb��Z�n�K�)��F�$� 11*ku[�FhJ��S�mY��to��p����^��/����z$Ί�?p^;�+���(��/X\��Mjo&I���V��W�%lAbI����W�j>����{B}to�g���zT@yh#C�e&L�Y�Q �GHp����܇'
e�Gs`��Ϭ ��bw�1������:�ڨ�IX��7)ۇ'� ��<uɃ��]�4�(=��;U:��ww>E<T�PA}� �	�t��U�Ȅ��?�U/ �Oׅ�RQ!�Vg~f.L��W�gO�Z��Ge�Ow�,�1�����6e0ό���p���$+_������|��;m����nc��&���p�����Γ�gx���>�g�S�꡸���Z�������mS����7��|9k��ڈ���w��,r�����ah�/4�ҡe��E�	�$�EDZ��La���1�dm�~��	�gd\�.^��Z)ǧ2�������[���~���o�'q�+�����.���
V�@�H�� ��@�N��);�0x�L"��oN��;���_j>AK��ͻ�Y����6-��:��.�=N1h2<.| ���?�7�����^�'k�I��!��WfO��,r�QJ,_�1Km�!���'�xb^��M�Z�Y��X�D��}b�1{;��n!j�O^^�Y�:+ �3e-���P���1խ��J�r8�$n��AC~�t�!�).�7"���\`�Q�0��<Y;g��������Ys�U�u�q��.�X;��a�q�2{�'���c�T�̅�<j����[L��v�)J���~��S��@ں �x��L��ضar��T'k����}-6��,��� �S�\�d7r��r�HJl�c�{Ӧ#�7Ĉ�x��./���э��LP��\��^bI)���\e�uN}A�.��r4+)4����Gv&��v�R=%vVk�*޳��$`�o�3��2�d8ۥG��\�͎q���!l:Yy*����?���F�y��{_<�Hv)��Eh���8�����h,A����K��J�	m�U|�FO��	l��&��k�A�A���Ś��L�7��QҞC���&K@�˕~���Xt\j6�eǓ��t:��NV d���<��ly�EG���9���׹�$4%�QA?7��P��ٯ�\g��&�z���3��ҿ�܄��x@�1�f6%0�76�����䭀T�g˂��矝�J=W� ���2�}*�Զ-k�݃Q�s	���59ш'l�� @E;B������/F���X�'���;D���>?-҆�:]�l%��3Gb��!��l< V^/�oe��Ȯ�O��>��Հ6#��\����'bj,�r/�q��9�}�^f�2޻��gf�n/�O)F4�X�%��-\�{�}��`������-��KN���K�U�1a8A��f�ӪK�x���4�T�&�K�� &�E�O/1���Gn��9}B����Ɨ0´�o�����{%�s���(+��^���O�=�RY�ӯj���a���FZ��l"sƴ-ޠ�2�rm��s�L�P�uk��� 0��~O�H+�~�����t��.��,!t��B�.N-u�I\I���t��#��!�@I���'Is��8�I��bB�7f���> ��e�WF=��Od��!�b�_)�����Is�n6�-�H��,r��yq78���|�����#��v�>cg���̯� o��a|3��p�:z��:-���4C߃Tqd����v��w=�l�܋�����Q`�ƫG�C�?����	m���2u9�_��&���ۿ�ebn��:���j18"�i�Uw:x�������3�	��x�
�{��. 3��-e����mEq�M6�f8��e�	�Y�����^�߸�Â�8�X����&�P8�.G�{�BM�}�u�xRO�V�#�7	�Z�-H�?������䝑-�������)l�(�~Y����d&�\+G�)��ݺ+�?M��,�׵�u(��ݾ�`]�O��0JW�G	���g�a|���-9�!��1㒝[���"��J����ؼ�N3{F����P�L��kⵜ���W��:B货4Im�2!��"�H����+��<�@\�>Al�uͮ��N���,�)k�d�Ώ�B��~d-5F�-
*�C���* �찢ꦻ��_T�F��]E_s^m�z��<k	�ě�\c��
O�(<�L:���G^��φ�+�/ ��ëk�tW�_�q��+�R3^0��Ul�$��d�Z�$�@Ѣ5]�o�����aj�%�\�~��h��a���%����h\�6��=m3�.w�TO�1q�Yõc�N�n�z.��9����l���W�S�gqK�*-�F�c��P�S4ts�%'�£5���g�F��j�f�5bf5Mhr�O��]s���,��� �Ѳ�3��-��YEH���	p�J�R�iApe[��<�<[����e��ʍe���6	M���8�u+Z�ޘ��%oQQ�y�筪	�?L1���QB;uBYA�Id�dC3R���@�������H���G-3@�]���T����.�_+�t���{��ki�?E��)y����*�3��S[>�W��`�c��g�|��n�T�j�D�Q�5C�򛄢��@��A�=���CN��v��- -���{��pN�$��zi�υ����t�?]Iǻ"��EE��sC+�O�M�"��]]�r���h=~���K �"�7wv�[��ݸ��s���'vø�L�J?�g�����z�"��Nߗ��u����?��
�%1'`n+�4�.�=L��s�SȞ&U�يT�Q�B��q�p���������e�T�xSߛУ+?<���(>�=�֐����8�G��w�`<��	SȽFY��g�讌��hL֗� h��6ˆf��#��*;�b��VFP	#HmDMw�Yu����H��b��A�A�F�G�*��+O��
-X�����������ʺ���`���,R���_�(���lv+G�R��/Hp�uK�۸&N��1��{^��l��F�dgP��~뻾�_�3���>5���}ҽ=@��U��r|�)QHA3�Z����+��T�L��n�*�$/\��d���8~��+�H��Yѐ��gopR�M��y��o[�8�&���8�cp7�^%�[q�lK�T�[,����yz9&&�Z�S��
��D�'�^���.W��i�A�o��8MY�m|Vn^o���e��d����+�~�C�Nj¢
��r��-sy��w��;T'�ү��Ȑ�	ء�#F�wV3{{��(??�7�`4]�N.n�pp䴗�7 �q�]	��A��uܸ��0ƿ���ѣ� �2b�5�G�Yj�i�j��ͩ���"Jwi��=	?X�U|�K��[�Gq��E�M�j�yj�[#k3B�GtC2�Ě�r���g�c�O�ء���AP��R�U�A���2�Kgc�������3;`��P��w��^7�S/����aI�Z�K�������L��@�"�==����*��G�@�>$�l���>��uļ��^1�7ϷU�������-�|��2��CAq3��#q&����ӡP>�Hs�vB!�l�@��x�!Ֆm/t���2-xX��f���۫E���<�l�/C{[C�tM���m��fK�/����',u���^�Bѩ�H�.
�I�cy����Q���CI�Z�&2i�Dq��l�&��ݾ��I�`]ܥz��`��aN|n�kr6��~���yG��/N%���M��HE�m}��!�j&^�jnZލ�ݷx��)Z$*�:�.d��ap���u.��z�^�Ɇ�ˑ�F�ܹ�,Vv;+�fG��]�&��{ӊ��܌
_�'�ats��9�J��_²��^����3���ԣ��������WK�M�����Q����Ň01�}���<���T�.w�튀�
2����)0�e��-��@=�.��H���?�.�j�hw^��:,��:z�ږƊ|n��*'�[s�r���c���9ٵZ��f`��jU�r 2���ĻVw�]��Z>-x��x=���V���(�%�_LfF���l�g0�z�̡C��8'5V3�Lu�f��GvRm�͔2z4�[^D��4
�-.b�Y�\�P���la�1�JY��50壈�&��S��v�!�4�O�cg��>���M���z�#��d���s�
�%���5��(!��5 R3-S��%��I�3��
hH���u�`����+�$��N��>���HW�s��d���F1���5���ƵǝCS�#g��~�೉I���*k[
�˵$� �tzj�h*��PE�m���'e�R�)_c��Oe����܍ "����2���(����z���O�ɥ�_'��A��+������~��=Z��������O��䧪/��f���
��ԩi����u@�'H��EI��`+�q����8+`Sa,!,H��u��Z�ZU�U�>-���wr=�\n��gM�*r�~v�_���Y!������9�9E���Є�_?17xV��`�N���YD�<���]=���:*Œf��=�V͹���QyD�F	_����H���P���j+p�sM����*����,`BAh��]��r�����c��C{Uvo�I����سB 
�%�v�截�i2�[PU�/�Z��z'K5�?��T�i2��.E���1�/�����-@�2�maH����E�Dك��X�''HB�`n�x��Yw�VV*�)/{�<�AS�_	�N�q�:	t4�g���)O&U�+��7�[]���xB ��`���\�@+� ��^�	��ˮX9�τjW��8nA7�t>��ʆ[Z�?��uV,`lO��f	>Gy�vU-{3JWW�#S:�I���� �� �1����GIm�_QRф).�iv{��h�ϫ��|HN�m���A[��AJa"G!����SlV�����==�"��Pt4Um~�+����y� ;�>�K���_l���6�3w��h�r�{�@a��a���C�)����P����=$�~t�1�Y�Ҁ��N�dr�vx�p��@����I>���p����u�Q��p�g�Ȗ�����i�K�ط����7ݿ+^/fD�6 ��M�M�8/�P�>T�@ad��$���P����::K�S�CN��TBD�y@��]C�D,��\����'��E_z��# ���8�W������;	�pbh��������+�Fd�sq{�:��S���PK   0jSU��Bv�  b     jsons/user_defined.json��ko�0��J���Q|w�m[��C �	%���$��4M��ػ��u��o�}�sl���o��V�,�[�|/�6�*�(����T�H�$��K��njξ�>��eW.���Re�57���yp�w���B�ujQ576"�l������q)�J2�@�dH�
�"����(��&�r\i������S1s�����}��"?鉏�W���U8���jn�z��UK���p����X]ߍ��1��ߛ�4�z[By\|�S.�&�	Uk\��f�"m(G��@��!n�����Uc����r�Ύ�U�2�x7]g��o���x4����wM՗��x���N�z���d�!�+Ww�}~��k�(���n�Z5��S��pY�#������N�N^��e*@�0$!9�� �9CL1�u:AX>���	K���'`1N¯(+�>EUd,}����c5%�I����;p(��>�Y�T򧏖P�0ʴRMl��&�r*�L'L<AK>x-��R{����}x��)�mW���bbp�Y�8>�*�<l�Ӄ��4��s�0]��Oj�.;���U�>}�"��%`i@B G�J���$��|B��=���FB4��ET�s(v�u�X��lb?��������h*|h�k8�
�/����Kg�蓏�o�O>S��>�P�mt�S��F2��/�Ue�dW5>���Bp�0�@�h$��cp�y���95�}�q]�4�-��}=[7�X���{|5G�;ѓ{�{_W�?PK
   0jSU:e!��&  �>                  cirkitFile.jsonPK
   �dSUv_Xh   t   /             '  images/0cd87e23-7b82-4f28-8831-3bf70f36678e.pngPK
   �]SUs� ^  7_  /             �'  images/12e44cfc-662f-4e22-b257-55fcd330266b.jpgPK
   |aSU��|�`  �c  /             �  images/290656fc-115e-450b-8d33-ab580af06883.jpgPK
   �[SU;��I�Y  \  /             ��  images/7842ad2d-d233-404b-8e7b-b5b626e67ff9.jpgPK
   �[SU;��I�Y  \  /             �@ images/943ec6f2-96cb-4ded-92cf-fc08d4cf4108.jpgPK
   0jSU��Bv�  b               � jsons/user_defined.jsonPK      S  �   